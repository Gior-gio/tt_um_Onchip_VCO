VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_Onchip_VCOx2
  CLASS BLOCK ;
  FOREIGN tt_um_Onchip_VCOx2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNADIFFAREA 1.800000 ;
    PORT
      LAYER li1 ;
        RECT 134.905 21.690 135.075 23.460 ;
        RECT 135.805 21.690 135.975 23.460 ;
        RECT 134.905 18.490 135.075 19.180 ;
        RECT 135.805 18.490 135.975 19.180 ;
      LAYER met1 ;
        RECT 134.875 21.960 135.105 23.440 ;
        RECT 135.775 21.960 136.005 23.440 ;
        RECT 134.825 21.690 135.155 21.960 ;
        RECT 135.725 21.690 136.055 21.960 ;
        RECT 136.945 21.480 137.745 21.510 ;
        RECT 134.825 21.210 137.745 21.480 ;
        RECT 136.945 21.180 137.745 21.210 ;
        RECT 134.875 19.145 135.105 19.160 ;
        RECT 135.775 19.145 136.005 19.160 ;
        RECT 134.830 18.885 135.150 19.145 ;
        RECT 135.730 18.885 136.050 19.145 ;
        RECT 134.875 18.510 135.105 18.885 ;
        RECT 135.775 18.510 136.005 18.885 ;
      LAYER met2 ;
        RECT 134.825 21.690 135.155 21.960 ;
        RECT 135.725 21.690 136.055 21.960 ;
        RECT 134.890 21.480 135.090 21.690 ;
        RECT 135.790 21.480 135.990 21.690 ;
        RECT 134.825 21.210 135.155 21.480 ;
        RECT 135.725 21.210 136.055 21.480 ;
        RECT 134.890 19.145 135.090 21.210 ;
        RECT 135.790 19.145 135.990 21.210 ;
        RECT 136.945 21.180 137.745 21.510 ;
        RECT 134.830 18.885 135.150 19.145 ;
        RECT 135.730 18.885 136.050 19.145 ;
      LAYER met3 ;
        RECT 136.945 21.180 152.710 21.510 ;
      LAYER met4 ;
        RECT 151.810 0.000 152.710 21.510 ;
    END
  END ua[0]
  PIN ua[2]
    ANTENNAGATEAREA 2.100000 ;
    PORT
      LAYER li1 ;
        RECT 127.170 19.535 127.520 19.805 ;
        RECT 131.070 19.535 131.420 19.805 ;
        RECT 123.920 11.325 124.270 11.595 ;
        RECT 125.870 11.325 126.220 11.595 ;
        RECT 129.770 11.325 130.120 11.595 ;
        RECT 133.670 11.325 134.020 11.595 ;
      LAYER met1 ;
        RECT 120.910 19.535 136.605 19.805 ;
        RECT 120.885 16.695 121.255 17.025 ;
        RECT 120.455 11.325 136.605 11.595 ;
      LAYER met2 ;
        RECT 120.910 19.535 121.230 19.805 ;
        RECT 120.935 17.025 121.205 19.535 ;
        RECT 120.885 16.695 121.255 17.025 ;
        RECT 120.935 11.595 121.205 16.695 ;
        RECT 120.910 11.325 121.230 11.595 ;
      LAYER met3 ;
        RECT 113.170 16.695 121.255 17.025 ;
      LAYER met4 ;
        RECT 113.170 0.000 114.070 17.025 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 1.800000 ;
    PORT
      LAYER li1 ;
        RECT 76.945 21.690 77.115 23.460 ;
        RECT 77.845 21.690 78.015 23.460 ;
        RECT 76.945 18.490 77.115 19.180 ;
        RECT 77.845 18.490 78.015 19.180 ;
      LAYER met1 ;
        RECT 76.915 21.960 77.145 23.440 ;
        RECT 77.815 21.960 78.045 23.440 ;
        RECT 76.865 21.690 77.195 21.960 ;
        RECT 77.765 21.690 78.095 21.960 ;
        RECT 78.985 21.480 79.785 21.510 ;
        RECT 76.865 21.210 79.785 21.480 ;
        RECT 78.985 21.180 79.785 21.210 ;
        RECT 76.915 19.145 77.145 19.160 ;
        RECT 77.815 19.145 78.045 19.160 ;
        RECT 76.870 18.885 77.190 19.145 ;
        RECT 77.770 18.885 78.090 19.145 ;
        RECT 76.915 18.510 77.145 18.885 ;
        RECT 77.815 18.510 78.045 18.885 ;
      LAYER met2 ;
        RECT 76.865 21.690 77.195 21.960 ;
        RECT 77.765 21.690 78.095 21.960 ;
        RECT 76.930 21.480 77.130 21.690 ;
        RECT 77.830 21.480 78.030 21.690 ;
        RECT 76.865 21.210 77.195 21.480 ;
        RECT 77.765 21.210 78.095 21.480 ;
        RECT 76.930 19.145 77.130 21.210 ;
        RECT 77.830 19.145 78.030 21.210 ;
        RECT 78.985 21.180 79.785 21.510 ;
        RECT 76.870 18.885 77.190 19.145 ;
        RECT 77.770 18.885 78.090 19.145 ;
      LAYER met3 ;
        RECT 78.985 21.180 94.750 21.510 ;
      LAYER met4 ;
        RECT 93.850 0.000 94.750 21.510 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNAGATEAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 64.980 16.065 65.310 16.395 ;
        RECT 66.620 16.145 66.950 16.315 ;
        RECT 68.570 16.145 68.900 16.315 ;
        RECT 70.520 16.145 70.850 16.315 ;
        RECT 72.470 16.145 72.800 16.315 ;
        RECT 74.420 16.145 74.750 16.315 ;
        RECT 66.620 14.815 66.950 14.985 ;
        RECT 68.570 14.815 68.900 14.985 ;
        RECT 70.520 14.815 70.850 14.985 ;
        RECT 72.470 14.815 72.800 14.985 ;
        RECT 74.420 14.815 74.750 14.985 ;
        RECT 76.370 14.815 76.700 14.985 ;
      LAYER met1 ;
        RECT 63.385 16.065 63.755 16.395 ;
        RECT 64.960 16.065 65.330 16.395 ;
        RECT 66.600 16.065 66.970 16.395 ;
        RECT 68.550 16.065 68.920 16.395 ;
        RECT 70.500 16.065 70.870 16.395 ;
        RECT 72.450 16.065 72.820 16.395 ;
        RECT 74.400 16.065 74.770 16.395 ;
        RECT 63.385 14.735 63.755 15.065 ;
        RECT 66.600 14.735 66.970 15.065 ;
        RECT 68.550 14.735 68.920 15.065 ;
        RECT 70.500 14.735 70.870 15.065 ;
        RECT 72.450 14.735 72.820 15.065 ;
        RECT 74.400 14.735 74.770 15.065 ;
        RECT 76.350 14.735 76.720 15.065 ;
      LAYER met2 ;
        RECT 63.385 16.065 63.755 16.395 ;
        RECT 64.960 16.065 65.330 16.395 ;
        RECT 66.600 16.065 66.970 16.395 ;
        RECT 68.550 16.065 68.920 16.395 ;
        RECT 70.500 16.065 70.870 16.395 ;
        RECT 72.450 16.065 72.820 16.395 ;
        RECT 74.400 16.065 74.770 16.395 ;
        RECT 63.435 15.065 63.705 16.065 ;
        RECT 63.385 14.735 63.755 15.065 ;
        RECT 66.600 14.735 66.970 15.065 ;
        RECT 68.550 14.735 68.920 15.065 ;
        RECT 70.500 14.735 70.870 15.065 ;
        RECT 72.450 14.735 72.820 15.065 ;
        RECT 74.400 14.735 74.770 15.065 ;
        RECT 76.350 14.735 76.720 15.065 ;
      LAYER met3 ;
        RECT 62.515 16.065 81.790 16.395 ;
        RECT 80.890 15.065 81.790 16.065 ;
        RECT 63.385 14.735 81.790 15.065 ;
      LAYER met4 ;
        RECT 80.890 2.400 81.790 16.395 ;
        RECT 74.530 1.500 81.790 2.400 ;
        RECT 74.530 0.000 75.430 1.500 ;
    END
  END ua[4]
  PIN ua[5]
    ANTENNAGATEAREA 2.100000 ;
    PORT
      LAYER li1 ;
        RECT 69.210 19.535 69.560 19.805 ;
        RECT 73.110 19.535 73.460 19.805 ;
        RECT 65.960 11.325 66.310 11.595 ;
        RECT 67.910 11.325 68.260 11.595 ;
        RECT 71.810 11.325 72.160 11.595 ;
        RECT 75.710 11.325 76.060 11.595 ;
      LAYER met1 ;
        RECT 62.950 19.535 78.645 19.805 ;
        RECT 62.925 16.695 63.295 17.025 ;
        RECT 62.495 11.325 78.645 11.595 ;
      LAYER met2 ;
        RECT 62.950 19.535 63.270 19.805 ;
        RECT 62.975 17.025 63.245 19.535 ;
        RECT 62.925 16.695 63.295 17.025 ;
        RECT 62.975 11.595 63.245 16.695 ;
        RECT 62.950 11.325 63.270 11.595 ;
      LAYER met3 ;
        RECT 55.210 16.695 63.295 17.025 ;
      LAYER met4 ;
        RECT 55.210 0.000 56.110 17.025 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNAGATEAREA 18.900000 ;
    ANTENNADIFFAREA 32.911999 ;
    PORT
      LAYER pwell ;
        RECT 66.180 18.205 78.210 19.465 ;
        RECT 124.140 18.205 136.170 19.465 ;
        RECT 66.180 17.725 77.765 18.205 ;
        RECT 124.140 17.725 135.725 18.205 ;
        RECT 64.880 17.535 77.765 17.725 ;
        RECT 122.840 17.535 135.725 17.725 ;
        RECT 64.880 15.895 75.840 17.535 ;
        RECT 122.840 15.895 133.800 17.535 ;
        RECT 64.860 15.235 77.640 15.895 ;
        RECT 122.820 15.235 135.600 15.895 ;
        RECT 65.530 14.665 77.640 15.235 ;
        RECT 123.490 14.665 135.600 15.235 ;
        RECT 65.530 13.405 77.790 14.665 ;
        RECT 123.490 13.405 135.750 14.665 ;
        RECT 65.530 11.665 77.140 13.405 ;
        RECT 123.490 11.665 135.100 13.405 ;
      LAYER li1 ;
        RECT 67.675 18.490 67.845 19.180 ;
        RECT 69.625 18.490 69.795 19.180 ;
        RECT 71.575 18.490 71.745 19.180 ;
        RECT 73.525 18.490 73.695 19.180 ;
        RECT 75.475 18.490 75.645 19.180 ;
        RECT 76.495 18.490 76.665 19.180 ;
        RECT 77.395 18.490 77.565 19.180 ;
        RECT 125.635 18.490 125.805 19.180 ;
        RECT 127.585 18.490 127.755 19.180 ;
        RECT 129.535 18.490 129.705 19.180 ;
        RECT 131.485 18.490 131.655 19.180 ;
        RECT 133.435 18.490 133.605 19.180 ;
        RECT 134.455 18.490 134.625 19.180 ;
        RECT 135.355 18.490 135.525 19.180 ;
        RECT 76.435 17.665 77.635 17.955 ;
        RECT 134.395 17.665 135.595 17.955 ;
        RECT 65.725 16.750 65.895 17.440 ;
        RECT 67.025 16.750 67.195 17.440 ;
        RECT 67.675 16.750 67.845 17.440 ;
        RECT 68.975 16.750 69.145 17.440 ;
        RECT 69.625 16.750 69.795 17.440 ;
        RECT 70.925 16.750 71.095 17.440 ;
        RECT 71.575 16.750 71.745 17.440 ;
        RECT 72.875 16.750 73.045 17.440 ;
        RECT 73.525 16.750 73.695 17.440 ;
        RECT 74.825 16.750 74.995 17.440 ;
        RECT 75.475 16.750 75.645 17.440 ;
        RECT 123.685 16.750 123.855 17.440 ;
        RECT 124.985 16.750 125.155 17.440 ;
        RECT 125.635 16.750 125.805 17.440 ;
        RECT 126.935 16.750 127.105 17.440 ;
        RECT 127.585 16.750 127.755 17.440 ;
        RECT 128.885 16.750 129.055 17.440 ;
        RECT 129.535 16.750 129.705 17.440 ;
        RECT 130.835 16.750 131.005 17.440 ;
        RECT 131.485 16.750 131.655 17.440 ;
        RECT 132.785 16.750 132.955 17.440 ;
        RECT 133.435 16.750 133.605 17.440 ;
        RECT 65.970 16.145 66.300 16.315 ;
        RECT 67.270 16.145 67.600 16.315 ;
        RECT 67.920 16.145 68.250 16.315 ;
        RECT 69.220 16.145 69.550 16.315 ;
        RECT 69.870 16.145 70.200 16.315 ;
        RECT 71.170 16.145 71.500 16.315 ;
        RECT 71.820 16.145 72.150 16.315 ;
        RECT 73.120 16.145 73.450 16.315 ;
        RECT 73.770 16.145 74.100 16.315 ;
        RECT 75.070 16.145 75.400 16.315 ;
        RECT 123.930 16.145 124.260 16.315 ;
        RECT 125.230 16.145 125.560 16.315 ;
        RECT 125.880 16.145 126.210 16.315 ;
        RECT 127.180 16.145 127.510 16.315 ;
        RECT 127.830 16.145 128.160 16.315 ;
        RECT 129.130 16.145 129.460 16.315 ;
        RECT 129.780 16.145 130.110 16.315 ;
        RECT 131.080 16.145 131.410 16.315 ;
        RECT 131.730 16.145 132.060 16.315 ;
        RECT 133.030 16.145 133.360 16.315 ;
        RECT 64.990 15.365 77.510 15.765 ;
        RECT 122.950 15.365 135.470 15.765 ;
        RECT 65.970 14.815 66.300 14.985 ;
        RECT 67.270 14.815 67.600 14.985 ;
        RECT 67.920 14.815 68.250 14.985 ;
        RECT 69.220 14.815 69.550 14.985 ;
        RECT 69.870 14.815 70.200 14.985 ;
        RECT 71.170 14.815 71.500 14.985 ;
        RECT 71.820 14.815 72.150 14.985 ;
        RECT 73.120 14.815 73.450 14.985 ;
        RECT 73.770 14.815 74.100 14.985 ;
        RECT 75.070 14.815 75.400 14.985 ;
        RECT 75.720 14.815 76.050 14.985 ;
        RECT 77.020 14.815 77.350 14.985 ;
        RECT 123.930 14.815 124.260 14.985 ;
        RECT 125.230 14.815 125.560 14.985 ;
        RECT 125.880 14.815 126.210 14.985 ;
        RECT 127.180 14.815 127.510 14.985 ;
        RECT 127.830 14.815 128.160 14.985 ;
        RECT 129.130 14.815 129.460 14.985 ;
        RECT 129.780 14.815 130.110 14.985 ;
        RECT 131.080 14.815 131.410 14.985 ;
        RECT 131.730 14.815 132.060 14.985 ;
        RECT 133.030 14.815 133.360 14.985 ;
        RECT 133.680 14.815 134.010 14.985 ;
        RECT 134.980 14.815 135.310 14.985 ;
        RECT 65.725 13.690 65.895 14.380 ;
        RECT 66.375 13.690 66.545 14.380 ;
        RECT 67.675 13.690 67.845 14.380 ;
        RECT 68.325 13.690 68.495 14.380 ;
        RECT 69.625 13.690 69.795 14.380 ;
        RECT 70.275 13.690 70.445 14.380 ;
        RECT 71.575 13.690 71.745 14.380 ;
        RECT 72.225 13.690 72.395 14.380 ;
        RECT 73.525 13.690 73.695 14.380 ;
        RECT 74.175 13.690 74.345 14.380 ;
        RECT 75.475 13.690 75.645 14.380 ;
        RECT 76.125 13.690 76.295 14.380 ;
        RECT 77.425 13.690 77.595 14.380 ;
        RECT 123.685 13.690 123.855 14.380 ;
        RECT 124.335 13.690 124.505 14.380 ;
        RECT 125.635 13.690 125.805 14.380 ;
        RECT 126.285 13.690 126.455 14.380 ;
        RECT 127.585 13.690 127.755 14.380 ;
        RECT 128.235 13.690 128.405 14.380 ;
        RECT 129.535 13.690 129.705 14.380 ;
        RECT 130.185 13.690 130.355 14.380 ;
        RECT 131.485 13.690 131.655 14.380 ;
        RECT 132.135 13.690 132.305 14.380 ;
        RECT 133.435 13.690 133.605 14.380 ;
        RECT 134.085 13.690 134.255 14.380 ;
        RECT 135.385 13.690 135.555 14.380 ;
        RECT 65.725 11.950 65.895 12.640 ;
        RECT 67.675 11.950 67.845 12.640 ;
        RECT 69.625 11.950 69.795 12.640 ;
        RECT 71.575 11.950 71.745 12.640 ;
        RECT 73.525 11.950 73.695 12.640 ;
        RECT 75.475 11.950 75.645 12.640 ;
        RECT 123.685 11.950 123.855 12.640 ;
        RECT 125.635 11.950 125.805 12.640 ;
        RECT 127.585 11.950 127.755 12.640 ;
        RECT 129.535 11.950 129.705 12.640 ;
        RECT 131.485 11.950 131.655 12.640 ;
        RECT 133.435 11.950 133.605 12.640 ;
      LAYER met1 ;
        RECT 67.600 18.510 67.920 19.160 ;
        RECT 69.550 18.510 69.870 19.160 ;
        RECT 71.500 18.510 71.820 19.160 ;
        RECT 73.450 18.510 73.770 19.160 ;
        RECT 75.400 18.510 75.720 19.160 ;
        RECT 76.465 18.785 76.695 19.160 ;
        RECT 77.365 18.785 77.595 19.160 ;
        RECT 76.420 18.525 76.740 18.785 ;
        RECT 77.320 18.525 77.640 18.785 ;
        RECT 76.465 18.510 76.695 18.525 ;
        RECT 77.365 18.510 77.595 18.525 ;
        RECT 125.560 18.510 125.880 19.160 ;
        RECT 127.510 18.510 127.830 19.160 ;
        RECT 129.460 18.510 129.780 19.160 ;
        RECT 131.410 18.510 131.730 19.160 ;
        RECT 133.360 18.510 133.680 19.160 ;
        RECT 134.425 18.785 134.655 19.160 ;
        RECT 135.325 18.785 135.555 19.160 ;
        RECT 134.380 18.525 134.700 18.785 ;
        RECT 135.280 18.525 135.600 18.785 ;
        RECT 134.425 18.510 134.655 18.525 ;
        RECT 135.325 18.510 135.555 18.525 ;
        RECT 76.435 17.665 77.635 17.955 ;
        RECT 134.395 17.665 135.595 17.955 ;
        RECT 65.695 17.345 65.925 17.420 ;
        RECT 66.995 17.345 67.225 17.420 ;
        RECT 67.645 17.345 67.875 17.420 ;
        RECT 68.945 17.345 69.175 17.420 ;
        RECT 69.595 17.345 69.825 17.420 ;
        RECT 70.895 17.345 71.125 17.420 ;
        RECT 71.545 17.345 71.775 17.420 ;
        RECT 72.845 17.345 73.075 17.420 ;
        RECT 73.495 17.345 73.725 17.420 ;
        RECT 74.795 17.345 75.025 17.420 ;
        RECT 75.445 17.345 75.675 17.420 ;
        RECT 123.655 17.345 123.885 17.420 ;
        RECT 124.955 17.345 125.185 17.420 ;
        RECT 125.605 17.345 125.835 17.420 ;
        RECT 126.905 17.345 127.135 17.420 ;
        RECT 127.555 17.345 127.785 17.420 ;
        RECT 128.855 17.345 129.085 17.420 ;
        RECT 129.505 17.345 129.735 17.420 ;
        RECT 130.805 17.345 131.035 17.420 ;
        RECT 131.455 17.345 131.685 17.420 ;
        RECT 132.755 17.345 132.985 17.420 ;
        RECT 133.405 17.345 133.635 17.420 ;
        RECT 65.625 16.845 65.995 17.345 ;
        RECT 66.925 16.845 67.295 17.345 ;
        RECT 67.575 16.845 67.945 17.345 ;
        RECT 68.875 16.845 69.245 17.345 ;
        RECT 69.525 16.845 69.895 17.345 ;
        RECT 70.825 16.845 71.195 17.345 ;
        RECT 71.475 16.845 71.845 17.345 ;
        RECT 72.775 16.845 73.145 17.345 ;
        RECT 73.425 16.845 73.795 17.345 ;
        RECT 74.725 16.845 75.095 17.345 ;
        RECT 75.375 16.845 75.745 17.345 ;
        RECT 123.585 16.845 123.955 17.345 ;
        RECT 124.885 16.845 125.255 17.345 ;
        RECT 125.535 16.845 125.905 17.345 ;
        RECT 126.835 16.845 127.205 17.345 ;
        RECT 127.485 16.845 127.855 17.345 ;
        RECT 128.785 16.845 129.155 17.345 ;
        RECT 129.435 16.845 129.805 17.345 ;
        RECT 130.735 16.845 131.105 17.345 ;
        RECT 131.385 16.845 131.755 17.345 ;
        RECT 132.685 16.845 133.055 17.345 ;
        RECT 133.335 16.845 133.705 17.345 ;
        RECT 65.695 16.770 65.925 16.845 ;
        RECT 66.995 16.770 67.225 16.845 ;
        RECT 67.645 16.770 67.875 16.845 ;
        RECT 68.945 16.770 69.175 16.845 ;
        RECT 69.595 16.770 69.825 16.845 ;
        RECT 70.895 16.770 71.125 16.845 ;
        RECT 71.545 16.770 71.775 16.845 ;
        RECT 72.845 16.770 73.075 16.845 ;
        RECT 73.495 16.770 73.725 16.845 ;
        RECT 74.795 16.770 75.025 16.845 ;
        RECT 75.445 16.770 75.675 16.845 ;
        RECT 123.655 16.770 123.885 16.845 ;
        RECT 124.955 16.770 125.185 16.845 ;
        RECT 125.605 16.770 125.835 16.845 ;
        RECT 126.905 16.770 127.135 16.845 ;
        RECT 127.555 16.770 127.785 16.845 ;
        RECT 128.855 16.770 129.085 16.845 ;
        RECT 129.505 16.770 129.735 16.845 ;
        RECT 130.805 16.770 131.035 16.845 ;
        RECT 131.455 16.770 131.685 16.845 ;
        RECT 132.755 16.770 132.985 16.845 ;
        RECT 133.405 16.770 133.635 16.845 ;
        RECT 65.950 15.765 66.320 16.345 ;
        RECT 67.250 15.765 67.620 16.345 ;
        RECT 67.900 15.765 68.270 16.345 ;
        RECT 69.200 15.765 69.570 16.345 ;
        RECT 69.850 15.765 70.220 16.345 ;
        RECT 71.150 15.765 71.520 16.345 ;
        RECT 71.800 15.765 72.170 16.345 ;
        RECT 73.100 15.765 73.470 16.345 ;
        RECT 73.750 15.765 74.120 16.345 ;
        RECT 75.050 15.765 75.420 16.345 ;
        RECT 123.910 15.765 124.280 16.345 ;
        RECT 125.210 15.765 125.580 16.345 ;
        RECT 125.860 15.765 126.230 16.345 ;
        RECT 127.160 15.765 127.530 16.345 ;
        RECT 127.810 15.765 128.180 16.345 ;
        RECT 129.110 15.765 129.480 16.345 ;
        RECT 129.760 15.765 130.130 16.345 ;
        RECT 131.060 15.765 131.430 16.345 ;
        RECT 131.710 15.765 132.080 16.345 ;
        RECT 133.010 15.765 133.380 16.345 ;
        RECT 64.990 15.365 77.510 15.765 ;
        RECT 122.950 15.365 135.470 15.765 ;
        RECT 65.950 14.785 66.320 15.365 ;
        RECT 67.250 14.785 67.620 15.365 ;
        RECT 67.900 14.785 68.270 15.365 ;
        RECT 69.200 14.785 69.570 15.365 ;
        RECT 69.850 14.785 70.220 15.365 ;
        RECT 71.150 14.785 71.520 15.365 ;
        RECT 71.800 14.785 72.170 15.365 ;
        RECT 73.100 14.785 73.470 15.365 ;
        RECT 73.750 14.785 74.120 15.365 ;
        RECT 75.050 14.785 75.420 15.365 ;
        RECT 75.700 14.785 76.070 15.365 ;
        RECT 77.000 14.785 77.370 15.365 ;
        RECT 123.910 14.785 124.280 15.365 ;
        RECT 125.210 14.785 125.580 15.365 ;
        RECT 125.860 14.785 126.230 15.365 ;
        RECT 127.160 14.785 127.530 15.365 ;
        RECT 127.810 14.785 128.180 15.365 ;
        RECT 129.110 14.785 129.480 15.365 ;
        RECT 129.760 14.785 130.130 15.365 ;
        RECT 131.060 14.785 131.430 15.365 ;
        RECT 131.710 14.785 132.080 15.365 ;
        RECT 133.010 14.785 133.380 15.365 ;
        RECT 133.660 14.785 134.030 15.365 ;
        RECT 134.960 14.785 135.330 15.365 ;
        RECT 65.695 14.285 65.925 14.360 ;
        RECT 66.345 14.285 66.575 14.360 ;
        RECT 67.645 14.285 67.875 14.360 ;
        RECT 68.295 14.285 68.525 14.360 ;
        RECT 69.595 14.285 69.825 14.360 ;
        RECT 70.245 14.285 70.475 14.360 ;
        RECT 71.545 14.285 71.775 14.360 ;
        RECT 72.195 14.285 72.425 14.360 ;
        RECT 73.495 14.285 73.725 14.360 ;
        RECT 74.145 14.285 74.375 14.360 ;
        RECT 75.445 14.285 75.675 14.360 ;
        RECT 76.095 14.285 76.325 14.360 ;
        RECT 77.395 14.285 77.625 14.360 ;
        RECT 123.655 14.285 123.885 14.360 ;
        RECT 124.305 14.285 124.535 14.360 ;
        RECT 125.605 14.285 125.835 14.360 ;
        RECT 126.255 14.285 126.485 14.360 ;
        RECT 127.555 14.285 127.785 14.360 ;
        RECT 128.205 14.285 128.435 14.360 ;
        RECT 129.505 14.285 129.735 14.360 ;
        RECT 130.155 14.285 130.385 14.360 ;
        RECT 131.455 14.285 131.685 14.360 ;
        RECT 132.105 14.285 132.335 14.360 ;
        RECT 133.405 14.285 133.635 14.360 ;
        RECT 134.055 14.285 134.285 14.360 ;
        RECT 135.355 14.285 135.585 14.360 ;
        RECT 65.625 13.785 65.995 14.285 ;
        RECT 66.275 13.785 66.645 14.285 ;
        RECT 67.575 13.785 67.945 14.285 ;
        RECT 68.225 13.785 68.595 14.285 ;
        RECT 69.525 13.785 69.895 14.285 ;
        RECT 70.175 13.785 70.545 14.285 ;
        RECT 71.475 13.785 71.845 14.285 ;
        RECT 72.125 13.785 72.495 14.285 ;
        RECT 73.425 13.785 73.795 14.285 ;
        RECT 74.075 13.785 74.445 14.285 ;
        RECT 75.375 13.785 75.745 14.285 ;
        RECT 76.025 13.785 76.395 14.285 ;
        RECT 77.325 13.785 77.695 14.285 ;
        RECT 123.585 13.785 123.955 14.285 ;
        RECT 124.235 13.785 124.605 14.285 ;
        RECT 125.535 13.785 125.905 14.285 ;
        RECT 126.185 13.785 126.555 14.285 ;
        RECT 127.485 13.785 127.855 14.285 ;
        RECT 128.135 13.785 128.505 14.285 ;
        RECT 129.435 13.785 129.805 14.285 ;
        RECT 130.085 13.785 130.455 14.285 ;
        RECT 131.385 13.785 131.755 14.285 ;
        RECT 132.035 13.785 132.405 14.285 ;
        RECT 133.335 13.785 133.705 14.285 ;
        RECT 133.985 13.785 134.355 14.285 ;
        RECT 135.285 13.785 135.655 14.285 ;
        RECT 65.695 13.710 65.925 13.785 ;
        RECT 66.345 13.710 66.575 13.785 ;
        RECT 67.645 13.710 67.875 13.785 ;
        RECT 68.295 13.710 68.525 13.785 ;
        RECT 69.595 13.710 69.825 13.785 ;
        RECT 70.245 13.710 70.475 13.785 ;
        RECT 71.545 13.710 71.775 13.785 ;
        RECT 72.195 13.710 72.425 13.785 ;
        RECT 73.495 13.710 73.725 13.785 ;
        RECT 74.145 13.710 74.375 13.785 ;
        RECT 75.445 13.710 75.675 13.785 ;
        RECT 76.095 13.710 76.325 13.785 ;
        RECT 77.395 13.710 77.625 13.785 ;
        RECT 123.655 13.710 123.885 13.785 ;
        RECT 124.305 13.710 124.535 13.785 ;
        RECT 125.605 13.710 125.835 13.785 ;
        RECT 126.255 13.710 126.485 13.785 ;
        RECT 127.555 13.710 127.785 13.785 ;
        RECT 128.205 13.710 128.435 13.785 ;
        RECT 129.505 13.710 129.735 13.785 ;
        RECT 130.155 13.710 130.385 13.785 ;
        RECT 131.455 13.710 131.685 13.785 ;
        RECT 132.105 13.710 132.335 13.785 ;
        RECT 133.405 13.710 133.635 13.785 ;
        RECT 134.055 13.710 134.285 13.785 ;
        RECT 135.355 13.710 135.585 13.785 ;
        RECT 65.650 11.970 65.970 12.620 ;
        RECT 67.600 11.970 67.920 12.620 ;
        RECT 69.550 11.970 69.870 12.620 ;
        RECT 71.500 11.970 71.820 12.620 ;
        RECT 73.450 11.970 73.770 12.620 ;
        RECT 75.400 11.970 75.720 12.620 ;
        RECT 123.610 11.970 123.930 12.620 ;
        RECT 125.560 11.970 125.880 12.620 ;
        RECT 127.510 11.970 127.830 12.620 ;
        RECT 129.460 11.970 129.780 12.620 ;
        RECT 131.410 11.970 131.730 12.620 ;
        RECT 133.360 11.970 133.680 12.620 ;
      LAYER met2 ;
        RECT 67.600 18.510 67.920 19.160 ;
        RECT 69.550 18.510 69.870 19.160 ;
        RECT 71.500 18.510 71.820 19.160 ;
        RECT 73.450 18.510 73.770 19.160 ;
        RECT 75.400 18.510 75.720 19.160 ;
        RECT 76.420 18.525 76.740 18.785 ;
        RECT 77.320 18.525 77.640 18.785 ;
        RECT 67.675 17.345 67.845 18.510 ;
        RECT 69.625 17.345 69.795 18.510 ;
        RECT 71.575 17.345 71.745 18.510 ;
        RECT 73.525 17.345 73.695 18.510 ;
        RECT 75.475 17.345 75.645 18.510 ;
        RECT 76.470 17.945 76.670 18.525 ;
        RECT 77.385 17.975 77.585 18.525 ;
        RECT 125.560 18.510 125.880 19.160 ;
        RECT 127.510 18.510 127.830 19.160 ;
        RECT 129.460 18.510 129.780 19.160 ;
        RECT 131.410 18.510 131.730 19.160 ;
        RECT 133.360 18.510 133.680 19.160 ;
        RECT 134.380 18.525 134.700 18.785 ;
        RECT 135.280 18.525 135.600 18.785 ;
        RECT 77.335 17.945 78.185 17.975 ;
        RECT 76.470 17.675 78.185 17.945 ;
        RECT 76.470 17.665 76.670 17.675 ;
        RECT 77.335 17.645 78.185 17.675 ;
        RECT 125.635 17.345 125.805 18.510 ;
        RECT 127.585 17.345 127.755 18.510 ;
        RECT 129.535 17.345 129.705 18.510 ;
        RECT 131.485 17.345 131.655 18.510 ;
        RECT 133.435 17.345 133.605 18.510 ;
        RECT 134.430 17.945 134.630 18.525 ;
        RECT 135.345 17.975 135.545 18.525 ;
        RECT 135.295 17.945 136.145 17.975 ;
        RECT 134.430 17.675 136.145 17.945 ;
        RECT 134.430 17.665 134.630 17.675 ;
        RECT 135.295 17.645 136.145 17.675 ;
        RECT 65.625 16.845 65.995 17.345 ;
        RECT 66.925 16.845 67.295 17.345 ;
        RECT 67.575 16.845 67.945 17.345 ;
        RECT 68.875 16.845 69.245 17.345 ;
        RECT 69.525 16.845 69.895 17.345 ;
        RECT 70.825 16.845 71.195 17.345 ;
        RECT 71.475 16.845 71.845 17.345 ;
        RECT 72.775 16.845 73.145 17.345 ;
        RECT 73.425 16.845 73.795 17.345 ;
        RECT 74.725 16.845 75.095 17.345 ;
        RECT 75.375 16.845 75.745 17.345 ;
        RECT 123.585 16.845 123.955 17.345 ;
        RECT 124.885 16.845 125.255 17.345 ;
        RECT 125.535 16.845 125.905 17.345 ;
        RECT 126.835 16.845 127.205 17.345 ;
        RECT 127.485 16.845 127.855 17.345 ;
        RECT 128.785 16.845 129.155 17.345 ;
        RECT 129.435 16.845 129.805 17.345 ;
        RECT 130.735 16.845 131.105 17.345 ;
        RECT 131.385 16.845 131.755 17.345 ;
        RECT 132.685 16.845 133.055 17.345 ;
        RECT 133.335 16.845 133.705 17.345 ;
        RECT 66.285 15.365 67.285 15.765 ;
        RECT 70.185 15.365 71.185 15.765 ;
        RECT 74.085 15.365 75.085 15.765 ;
        RECT 124.245 15.365 125.245 15.765 ;
        RECT 128.145 15.365 129.145 15.765 ;
        RECT 132.045 15.365 133.045 15.765 ;
        RECT 65.625 13.785 65.995 14.285 ;
        RECT 66.275 13.785 66.645 14.285 ;
        RECT 67.575 13.785 67.945 14.285 ;
        RECT 68.225 13.785 68.595 14.285 ;
        RECT 69.525 13.785 69.895 14.285 ;
        RECT 70.175 13.785 70.545 14.285 ;
        RECT 71.475 13.785 71.845 14.285 ;
        RECT 72.125 13.785 72.495 14.285 ;
        RECT 73.425 13.785 73.795 14.285 ;
        RECT 74.075 13.785 74.445 14.285 ;
        RECT 75.375 13.785 75.745 14.285 ;
        RECT 76.025 13.785 76.395 14.285 ;
        RECT 77.325 13.785 77.695 14.285 ;
        RECT 123.585 13.785 123.955 14.285 ;
        RECT 124.235 13.785 124.605 14.285 ;
        RECT 125.535 13.785 125.905 14.285 ;
        RECT 126.185 13.785 126.555 14.285 ;
        RECT 127.485 13.785 127.855 14.285 ;
        RECT 128.135 13.785 128.505 14.285 ;
        RECT 129.435 13.785 129.805 14.285 ;
        RECT 130.085 13.785 130.455 14.285 ;
        RECT 131.385 13.785 131.755 14.285 ;
        RECT 132.035 13.785 132.405 14.285 ;
        RECT 133.335 13.785 133.705 14.285 ;
        RECT 133.985 13.785 134.355 14.285 ;
        RECT 135.285 13.785 135.655 14.285 ;
        RECT 65.725 12.620 65.895 13.785 ;
        RECT 67.675 12.620 67.845 13.785 ;
        RECT 69.625 12.620 69.795 13.785 ;
        RECT 71.575 12.620 71.745 13.785 ;
        RECT 73.525 12.620 73.695 13.785 ;
        RECT 75.475 12.620 75.645 13.785 ;
        RECT 123.685 12.620 123.855 13.785 ;
        RECT 125.635 12.620 125.805 13.785 ;
        RECT 127.585 12.620 127.755 13.785 ;
        RECT 129.535 12.620 129.705 13.785 ;
        RECT 131.485 12.620 131.655 13.785 ;
        RECT 133.435 12.620 133.605 13.785 ;
        RECT 65.650 11.970 65.970 12.620 ;
        RECT 67.600 11.970 67.920 12.620 ;
        RECT 69.550 11.970 69.870 12.620 ;
        RECT 71.500 11.970 71.820 12.620 ;
        RECT 73.450 11.970 73.770 12.620 ;
        RECT 75.400 11.970 75.720 12.620 ;
        RECT 123.610 11.970 123.930 12.620 ;
        RECT 125.560 11.970 125.880 12.620 ;
        RECT 127.510 11.970 127.830 12.620 ;
        RECT 129.460 11.970 129.780 12.620 ;
        RECT 131.410 11.970 131.730 12.620 ;
        RECT 133.360 11.970 133.680 12.620 ;
      LAYER met3 ;
        RECT 1.000 30.595 136.945 32.595 ;
        RECT 77.335 17.645 78.185 17.975 ;
        RECT 135.295 17.645 136.145 17.975 ;
        RECT 64.115 16.845 78.645 17.345 ;
        RECT 122.075 16.845 136.605 17.345 ;
        RECT 66.285 15.365 67.285 15.765 ;
        RECT 70.185 15.365 71.185 15.765 ;
        RECT 74.085 15.365 75.085 15.765 ;
        RECT 124.245 15.365 125.245 15.765 ;
        RECT 128.145 15.365 129.145 15.765 ;
        RECT 132.045 15.365 133.045 15.765 ;
        RECT 65.625 13.785 77.695 14.285 ;
        RECT 123.585 13.785 135.655 14.285 ;
      LAYER met4 ;
        RECT 30.670 220.760 30.970 225.760 ;
        RECT 33.430 220.760 33.730 225.760 ;
        RECT 36.190 220.760 36.490 225.760 ;
        RECT 38.950 220.760 39.250 225.760 ;
        RECT 41.710 220.760 42.010 225.760 ;
        RECT 44.470 220.760 44.770 225.760 ;
        RECT 47.230 220.760 47.530 225.760 ;
        RECT 49.990 220.760 50.290 225.760 ;
        RECT 52.750 220.760 53.050 225.760 ;
        RECT 55.510 220.760 55.810 225.760 ;
        RECT 58.270 220.760 58.570 225.760 ;
        RECT 61.030 220.760 61.330 225.760 ;
        RECT 63.790 220.760 64.090 225.760 ;
        RECT 66.550 220.760 66.850 225.760 ;
        RECT 69.310 220.760 69.610 225.760 ;
        RECT 72.070 220.760 72.370 225.760 ;
        RECT 74.830 220.760 75.130 225.760 ;
        RECT 77.590 220.760 77.890 225.760 ;
        RECT 80.350 220.760 80.650 225.760 ;
        RECT 83.110 220.760 83.410 225.760 ;
        RECT 85.870 220.760 86.170 225.760 ;
        RECT 88.630 220.760 88.930 225.760 ;
        RECT 91.390 220.760 91.690 225.760 ;
        RECT 94.150 220.760 94.450 225.760 ;
        RECT 4.000 219.760 94.450 220.760 ;
        RECT 4.000 5.000 6.000 219.760 ;
        RECT 62.150 3.585 63.150 37.250 ;
        RECT 66.285 3.585 67.285 37.250 ;
        RECT 70.185 3.585 71.185 37.250 ;
        RECT 74.085 3.585 75.085 37.250 ;
        RECT 77.985 17.975 78.985 37.250 ;
        RECT 77.335 17.645 78.985 17.975 ;
        RECT 77.985 3.585 78.985 17.645 ;
        RECT 120.110 3.585 121.110 37.250 ;
        RECT 124.245 3.585 125.245 37.250 ;
        RECT 128.145 3.585 129.145 37.250 ;
        RECT 132.045 3.585 133.045 37.250 ;
        RECT 135.945 17.975 136.945 37.250 ;
        RECT 135.295 17.645 136.945 17.975 ;
        RECT 135.945 3.585 136.945 17.645 ;
    END
  END uio_oe[0]
  PIN VDPWR
    ANTENNAGATEAREA 30.799999 ;
    ANTENNADIFFAREA 49.711998 ;
    PORT
      LAYER nwell ;
        RECT 64.705 23.955 77.965 27.725 ;
        RECT 122.665 23.955 135.925 27.725 ;
        RECT 64.705 21.195 78.385 23.955 ;
        RECT 122.665 21.195 136.345 23.955 ;
        RECT 64.705 20.855 77.965 21.195 ;
        RECT 122.665 20.855 135.925 21.195 ;
        RECT 64.705 3.405 77.965 10.275 ;
        RECT 122.665 3.405 135.925 10.275 ;
      LAYER li1 ;
        RECT 64.990 27.145 75.560 27.545 ;
        RECT 122.950 27.145 133.520 27.545 ;
        RECT 65.970 26.595 66.300 26.765 ;
        RECT 67.270 26.595 67.600 26.765 ;
        RECT 67.920 26.595 68.250 26.765 ;
        RECT 69.220 26.595 69.550 26.765 ;
        RECT 69.870 26.595 70.200 26.765 ;
        RECT 71.170 26.595 71.500 26.765 ;
        RECT 71.820 26.595 72.150 26.765 ;
        RECT 73.120 26.595 73.450 26.765 ;
        RECT 73.770 26.595 74.100 26.765 ;
        RECT 75.070 26.595 75.400 26.765 ;
        RECT 123.930 26.595 124.260 26.765 ;
        RECT 125.230 26.595 125.560 26.765 ;
        RECT 125.880 26.595 126.210 26.765 ;
        RECT 127.180 26.595 127.510 26.765 ;
        RECT 127.830 26.595 128.160 26.765 ;
        RECT 129.130 26.595 129.460 26.765 ;
        RECT 129.780 26.595 130.110 26.765 ;
        RECT 131.080 26.595 131.410 26.765 ;
        RECT 131.730 26.595 132.060 26.765 ;
        RECT 133.030 26.595 133.360 26.765 ;
        RECT 65.725 24.430 65.895 26.200 ;
        RECT 67.025 24.430 67.195 26.200 ;
        RECT 67.675 24.430 67.845 26.200 ;
        RECT 68.975 24.430 69.145 26.200 ;
        RECT 69.625 24.430 69.795 26.200 ;
        RECT 70.925 24.430 71.095 26.200 ;
        RECT 71.575 24.430 71.745 26.200 ;
        RECT 72.875 24.430 73.045 26.200 ;
        RECT 73.525 24.430 73.695 26.200 ;
        RECT 74.825 24.430 74.995 26.200 ;
        RECT 75.475 24.430 75.645 26.200 ;
        RECT 76.420 24.345 77.620 24.635 ;
        RECT 123.685 24.430 123.855 26.200 ;
        RECT 124.985 24.430 125.155 26.200 ;
        RECT 125.635 24.430 125.805 26.200 ;
        RECT 126.935 24.430 127.105 26.200 ;
        RECT 127.585 24.430 127.755 26.200 ;
        RECT 128.885 24.430 129.055 26.200 ;
        RECT 129.535 24.430 129.705 26.200 ;
        RECT 130.835 24.430 131.005 26.200 ;
        RECT 131.485 24.430 131.655 26.200 ;
        RECT 132.785 24.430 132.955 26.200 ;
        RECT 133.435 24.430 133.605 26.200 ;
        RECT 134.380 24.345 135.580 24.635 ;
        RECT 76.495 21.690 76.665 23.460 ;
        RECT 77.395 21.690 77.565 23.460 ;
        RECT 134.455 21.690 134.625 23.460 ;
        RECT 135.355 21.690 135.525 23.460 ;
        RECT 65.725 4.930 65.895 6.700 ;
        RECT 66.375 4.930 66.545 6.700 ;
        RECT 67.675 4.930 67.845 6.700 ;
        RECT 68.325 4.930 68.495 6.700 ;
        RECT 69.625 4.930 69.795 6.700 ;
        RECT 70.275 4.930 70.445 6.700 ;
        RECT 71.575 4.930 71.745 6.700 ;
        RECT 72.225 4.930 72.395 6.700 ;
        RECT 73.525 4.930 73.695 6.700 ;
        RECT 74.175 4.930 74.345 6.700 ;
        RECT 75.475 4.930 75.645 6.700 ;
        RECT 76.125 4.930 76.295 6.700 ;
        RECT 77.425 4.930 77.595 6.700 ;
        RECT 123.685 4.930 123.855 6.700 ;
        RECT 124.335 4.930 124.505 6.700 ;
        RECT 125.635 4.930 125.805 6.700 ;
        RECT 126.285 4.930 126.455 6.700 ;
        RECT 127.585 4.930 127.755 6.700 ;
        RECT 128.235 4.930 128.405 6.700 ;
        RECT 129.535 4.930 129.705 6.700 ;
        RECT 130.185 4.930 130.355 6.700 ;
        RECT 131.485 4.930 131.655 6.700 ;
        RECT 132.135 4.930 132.305 6.700 ;
        RECT 133.435 4.930 133.605 6.700 ;
        RECT 134.085 4.930 134.255 6.700 ;
        RECT 135.385 4.930 135.555 6.700 ;
        RECT 65.970 4.365 66.300 4.535 ;
        RECT 67.270 4.365 67.600 4.535 ;
        RECT 67.920 4.365 68.250 4.535 ;
        RECT 69.220 4.365 69.550 4.535 ;
        RECT 69.870 4.365 70.200 4.535 ;
        RECT 71.170 4.365 71.500 4.535 ;
        RECT 71.820 4.365 72.150 4.535 ;
        RECT 73.120 4.365 73.450 4.535 ;
        RECT 73.770 4.365 74.100 4.535 ;
        RECT 75.070 4.365 75.400 4.535 ;
        RECT 75.720 4.365 76.050 4.535 ;
        RECT 77.020 4.365 77.350 4.535 ;
        RECT 123.930 4.365 124.260 4.535 ;
        RECT 125.230 4.365 125.560 4.535 ;
        RECT 125.880 4.365 126.210 4.535 ;
        RECT 127.180 4.365 127.510 4.535 ;
        RECT 127.830 4.365 128.160 4.535 ;
        RECT 129.130 4.365 129.460 4.535 ;
        RECT 129.780 4.365 130.110 4.535 ;
        RECT 131.080 4.365 131.410 4.535 ;
        RECT 131.730 4.365 132.060 4.535 ;
        RECT 133.030 4.365 133.360 4.535 ;
        RECT 133.680 4.365 134.010 4.535 ;
        RECT 134.980 4.365 135.310 4.535 ;
        RECT 65.810 3.585 77.510 3.985 ;
        RECT 123.770 3.585 135.470 3.985 ;
      LAYER met1 ;
        RECT 64.115 27.145 77.965 27.545 ;
        RECT 122.075 27.145 135.925 27.545 ;
        RECT 65.950 26.565 66.320 27.145 ;
        RECT 67.250 26.565 67.620 27.145 ;
        RECT 67.900 26.565 68.270 27.145 ;
        RECT 69.200 26.565 69.570 27.145 ;
        RECT 69.850 26.565 70.220 27.145 ;
        RECT 71.150 26.565 71.520 27.145 ;
        RECT 71.800 26.565 72.170 27.145 ;
        RECT 73.100 26.565 73.470 27.145 ;
        RECT 73.750 26.565 74.120 27.145 ;
        RECT 75.050 26.565 75.420 27.145 ;
        RECT 123.910 26.565 124.280 27.145 ;
        RECT 125.210 26.565 125.580 27.145 ;
        RECT 125.860 26.565 126.230 27.145 ;
        RECT 127.160 26.565 127.530 27.145 ;
        RECT 127.810 26.565 128.180 27.145 ;
        RECT 129.110 26.565 129.480 27.145 ;
        RECT 129.760 26.565 130.130 27.145 ;
        RECT 131.060 26.565 131.430 27.145 ;
        RECT 131.710 26.565 132.080 27.145 ;
        RECT 133.010 26.565 133.380 27.145 ;
        RECT 65.695 25.565 65.925 26.180 ;
        RECT 66.995 25.565 67.225 26.180 ;
        RECT 67.645 25.565 67.875 26.180 ;
        RECT 68.945 25.565 69.175 26.180 ;
        RECT 69.595 25.565 69.825 26.180 ;
        RECT 70.895 25.565 71.125 26.180 ;
        RECT 71.545 25.565 71.775 26.180 ;
        RECT 72.845 25.565 73.075 26.180 ;
        RECT 73.495 25.565 73.725 26.180 ;
        RECT 74.795 25.565 75.025 26.180 ;
        RECT 75.445 25.565 75.675 26.180 ;
        RECT 123.655 25.565 123.885 26.180 ;
        RECT 124.955 25.565 125.185 26.180 ;
        RECT 125.605 25.565 125.835 26.180 ;
        RECT 126.905 25.565 127.135 26.180 ;
        RECT 127.555 25.565 127.785 26.180 ;
        RECT 128.855 25.565 129.085 26.180 ;
        RECT 129.505 25.565 129.735 26.180 ;
        RECT 130.805 25.565 131.035 26.180 ;
        RECT 131.455 25.565 131.685 26.180 ;
        RECT 132.755 25.565 132.985 26.180 ;
        RECT 133.405 25.565 133.635 26.180 ;
        RECT 65.625 25.065 65.995 25.565 ;
        RECT 66.925 25.065 67.295 25.565 ;
        RECT 67.575 25.065 67.945 25.565 ;
        RECT 68.875 25.065 69.245 25.565 ;
        RECT 69.525 25.065 69.895 25.565 ;
        RECT 70.825 25.065 71.195 25.565 ;
        RECT 71.475 25.065 71.845 25.565 ;
        RECT 72.775 25.065 73.145 25.565 ;
        RECT 73.425 25.065 73.795 25.565 ;
        RECT 74.725 25.065 75.095 25.565 ;
        RECT 75.375 25.065 75.745 25.565 ;
        RECT 123.585 25.065 123.955 25.565 ;
        RECT 124.885 25.065 125.255 25.565 ;
        RECT 125.535 25.065 125.905 25.565 ;
        RECT 126.835 25.065 127.205 25.565 ;
        RECT 127.485 25.065 127.855 25.565 ;
        RECT 128.785 25.065 129.155 25.565 ;
        RECT 129.435 25.065 129.805 25.565 ;
        RECT 130.735 25.065 131.105 25.565 ;
        RECT 131.385 25.065 131.755 25.565 ;
        RECT 132.685 25.065 133.055 25.565 ;
        RECT 133.335 25.065 133.705 25.565 ;
        RECT 65.695 24.450 65.925 25.065 ;
        RECT 66.995 24.450 67.225 25.065 ;
        RECT 67.645 24.450 67.875 25.065 ;
        RECT 68.945 24.450 69.175 25.065 ;
        RECT 69.595 24.450 69.825 25.065 ;
        RECT 70.895 24.450 71.125 25.065 ;
        RECT 71.545 24.450 71.775 25.065 ;
        RECT 72.845 24.450 73.075 25.065 ;
        RECT 73.495 24.450 73.725 25.065 ;
        RECT 74.795 24.450 75.025 25.065 ;
        RECT 75.445 24.450 75.675 25.065 ;
        RECT 76.420 24.345 77.620 24.635 ;
        RECT 123.655 24.450 123.885 25.065 ;
        RECT 124.955 24.450 125.185 25.065 ;
        RECT 125.605 24.450 125.835 25.065 ;
        RECT 126.905 24.450 127.135 25.065 ;
        RECT 127.555 24.450 127.785 25.065 ;
        RECT 128.855 24.450 129.085 25.065 ;
        RECT 129.505 24.450 129.735 25.065 ;
        RECT 130.805 24.450 131.035 25.065 ;
        RECT 131.455 24.450 131.685 25.065 ;
        RECT 132.755 24.450 132.985 25.065 ;
        RECT 133.405 24.450 133.635 25.065 ;
        RECT 134.380 24.345 135.580 24.635 ;
        RECT 76.465 23.425 76.695 23.440 ;
        RECT 77.365 23.425 77.595 23.440 ;
        RECT 134.425 23.425 134.655 23.440 ;
        RECT 135.325 23.425 135.555 23.440 ;
        RECT 76.420 23.165 76.740 23.425 ;
        RECT 77.320 23.165 77.640 23.425 ;
        RECT 134.380 23.165 134.700 23.425 ;
        RECT 135.280 23.165 135.600 23.425 ;
        RECT 76.465 21.710 76.695 23.165 ;
        RECT 77.365 21.710 77.595 23.165 ;
        RECT 134.425 21.710 134.655 23.165 ;
        RECT 135.325 21.710 135.555 23.165 ;
        RECT 65.695 6.065 65.925 6.680 ;
        RECT 66.345 6.065 66.575 6.680 ;
        RECT 67.645 6.065 67.875 6.680 ;
        RECT 68.295 6.065 68.525 6.680 ;
        RECT 69.595 6.065 69.825 6.680 ;
        RECT 70.245 6.065 70.475 6.680 ;
        RECT 71.545 6.065 71.775 6.680 ;
        RECT 72.195 6.065 72.425 6.680 ;
        RECT 73.495 6.065 73.725 6.680 ;
        RECT 74.145 6.065 74.375 6.680 ;
        RECT 75.445 6.065 75.675 6.680 ;
        RECT 76.095 6.065 76.325 6.680 ;
        RECT 77.395 6.065 77.625 6.680 ;
        RECT 123.655 6.065 123.885 6.680 ;
        RECT 124.305 6.065 124.535 6.680 ;
        RECT 125.605 6.065 125.835 6.680 ;
        RECT 126.255 6.065 126.485 6.680 ;
        RECT 127.555 6.065 127.785 6.680 ;
        RECT 128.205 6.065 128.435 6.680 ;
        RECT 129.505 6.065 129.735 6.680 ;
        RECT 130.155 6.065 130.385 6.680 ;
        RECT 131.455 6.065 131.685 6.680 ;
        RECT 132.105 6.065 132.335 6.680 ;
        RECT 133.405 6.065 133.635 6.680 ;
        RECT 134.055 6.065 134.285 6.680 ;
        RECT 135.355 6.065 135.585 6.680 ;
        RECT 65.625 5.565 65.995 6.065 ;
        RECT 66.275 5.565 66.645 6.065 ;
        RECT 67.575 5.565 67.945 6.065 ;
        RECT 68.225 5.565 68.595 6.065 ;
        RECT 69.525 5.565 69.895 6.065 ;
        RECT 70.175 5.565 70.545 6.065 ;
        RECT 71.475 5.565 71.845 6.065 ;
        RECT 72.125 5.565 72.495 6.065 ;
        RECT 73.425 5.565 73.795 6.065 ;
        RECT 74.075 5.565 74.445 6.065 ;
        RECT 75.375 5.565 75.745 6.065 ;
        RECT 76.025 5.565 76.395 6.065 ;
        RECT 77.325 5.565 77.695 6.065 ;
        RECT 123.585 5.565 123.955 6.065 ;
        RECT 124.235 5.565 124.605 6.065 ;
        RECT 125.535 5.565 125.905 6.065 ;
        RECT 126.185 5.565 126.555 6.065 ;
        RECT 127.485 5.565 127.855 6.065 ;
        RECT 128.135 5.565 128.505 6.065 ;
        RECT 129.435 5.565 129.805 6.065 ;
        RECT 130.085 5.565 130.455 6.065 ;
        RECT 131.385 5.565 131.755 6.065 ;
        RECT 132.035 5.565 132.405 6.065 ;
        RECT 133.335 5.565 133.705 6.065 ;
        RECT 133.985 5.565 134.355 6.065 ;
        RECT 135.285 5.565 135.655 6.065 ;
        RECT 65.695 4.950 65.925 5.565 ;
        RECT 66.345 4.950 66.575 5.565 ;
        RECT 67.645 4.950 67.875 5.565 ;
        RECT 68.295 4.950 68.525 5.565 ;
        RECT 69.595 4.950 69.825 5.565 ;
        RECT 70.245 4.950 70.475 5.565 ;
        RECT 71.545 4.950 71.775 5.565 ;
        RECT 72.195 4.950 72.425 5.565 ;
        RECT 73.495 4.950 73.725 5.565 ;
        RECT 74.145 4.950 74.375 5.565 ;
        RECT 75.445 4.950 75.675 5.565 ;
        RECT 76.095 4.950 76.325 5.565 ;
        RECT 77.395 4.950 77.625 5.565 ;
        RECT 123.655 4.950 123.885 5.565 ;
        RECT 124.305 4.950 124.535 5.565 ;
        RECT 125.605 4.950 125.835 5.565 ;
        RECT 126.255 4.950 126.485 5.565 ;
        RECT 127.555 4.950 127.785 5.565 ;
        RECT 128.205 4.950 128.435 5.565 ;
        RECT 129.505 4.950 129.735 5.565 ;
        RECT 130.155 4.950 130.385 5.565 ;
        RECT 131.455 4.950 131.685 5.565 ;
        RECT 132.105 4.950 132.335 5.565 ;
        RECT 133.405 4.950 133.635 5.565 ;
        RECT 134.055 4.950 134.285 5.565 ;
        RECT 135.355 4.950 135.585 5.565 ;
        RECT 65.950 3.985 66.320 4.565 ;
        RECT 67.250 3.985 67.620 4.565 ;
        RECT 67.900 3.985 68.270 4.565 ;
        RECT 69.200 3.985 69.570 4.565 ;
        RECT 69.850 3.985 70.220 4.565 ;
        RECT 71.150 3.985 71.520 4.565 ;
        RECT 71.800 3.985 72.170 4.565 ;
        RECT 73.100 3.985 73.470 4.565 ;
        RECT 73.750 3.985 74.120 4.565 ;
        RECT 75.050 3.985 75.420 4.565 ;
        RECT 75.700 3.985 76.070 4.565 ;
        RECT 77.000 3.985 77.370 4.565 ;
        RECT 123.910 3.985 124.280 4.565 ;
        RECT 125.210 3.985 125.580 4.565 ;
        RECT 125.860 3.985 126.230 4.565 ;
        RECT 127.160 3.985 127.530 4.565 ;
        RECT 127.810 3.985 128.180 4.565 ;
        RECT 129.110 3.985 129.480 4.565 ;
        RECT 129.760 3.985 130.130 4.565 ;
        RECT 131.060 3.985 131.430 4.565 ;
        RECT 131.710 3.985 132.080 4.565 ;
        RECT 133.010 3.985 133.380 4.565 ;
        RECT 133.660 3.985 134.030 4.565 ;
        RECT 134.960 3.985 135.330 4.565 ;
        RECT 64.115 3.585 78.485 3.985 ;
        RECT 122.075 3.585 136.445 3.985 ;
      LAYER met2 ;
        RECT 64.115 27.145 65.115 27.545 ;
        RECT 68.235 27.145 69.235 27.545 ;
        RECT 72.135 27.145 73.135 27.545 ;
        RECT 76.035 27.145 77.035 27.545 ;
        RECT 122.075 27.145 123.075 27.545 ;
        RECT 126.195 27.145 127.195 27.545 ;
        RECT 130.095 27.145 131.095 27.545 ;
        RECT 133.995 27.145 134.995 27.545 ;
        RECT 65.625 25.065 65.995 25.565 ;
        RECT 66.925 25.065 67.295 25.565 ;
        RECT 67.575 25.065 67.945 25.565 ;
        RECT 68.875 25.065 69.245 25.565 ;
        RECT 69.525 25.065 69.895 25.565 ;
        RECT 70.825 25.065 71.195 25.565 ;
        RECT 71.475 25.065 71.845 25.565 ;
        RECT 72.775 25.065 73.145 25.565 ;
        RECT 73.425 25.065 73.795 25.565 ;
        RECT 74.725 25.065 75.095 25.565 ;
        RECT 75.375 25.065 75.745 25.565 ;
        RECT 123.585 25.065 123.955 25.565 ;
        RECT 124.885 25.065 125.255 25.565 ;
        RECT 125.535 25.065 125.905 25.565 ;
        RECT 126.835 25.065 127.205 25.565 ;
        RECT 127.485 25.065 127.855 25.565 ;
        RECT 128.785 25.065 129.155 25.565 ;
        RECT 129.435 25.065 129.805 25.565 ;
        RECT 130.735 25.065 131.105 25.565 ;
        RECT 131.385 25.065 131.755 25.565 ;
        RECT 132.685 25.065 133.055 25.565 ;
        RECT 133.335 25.065 133.705 25.565 ;
        RECT 76.035 24.625 77.035 24.655 ;
        RECT 133.995 24.625 134.995 24.655 ;
        RECT 76.035 24.355 77.590 24.625 ;
        RECT 133.995 24.355 135.550 24.625 ;
        RECT 76.035 24.325 77.035 24.355 ;
        RECT 76.490 23.425 76.690 24.325 ;
        RECT 77.375 23.425 77.575 24.355 ;
        RECT 133.995 24.325 134.995 24.355 ;
        RECT 134.450 23.425 134.650 24.325 ;
        RECT 135.335 23.425 135.535 24.355 ;
        RECT 76.420 23.165 76.740 23.425 ;
        RECT 77.320 23.165 77.640 23.425 ;
        RECT 134.380 23.165 134.700 23.425 ;
        RECT 135.280 23.165 135.600 23.425 ;
        RECT 65.625 5.565 65.995 6.065 ;
        RECT 66.275 5.565 66.645 6.065 ;
        RECT 67.575 5.565 67.945 6.065 ;
        RECT 68.225 5.565 68.595 6.065 ;
        RECT 69.525 5.565 69.895 6.065 ;
        RECT 70.175 5.565 70.545 6.065 ;
        RECT 71.475 5.565 71.845 6.065 ;
        RECT 72.125 5.565 72.495 6.065 ;
        RECT 73.425 5.565 73.795 6.065 ;
        RECT 74.075 5.565 74.445 6.065 ;
        RECT 75.375 5.565 75.745 6.065 ;
        RECT 76.025 5.565 76.395 6.065 ;
        RECT 77.325 5.565 77.695 6.065 ;
        RECT 123.585 5.565 123.955 6.065 ;
        RECT 124.235 5.565 124.605 6.065 ;
        RECT 125.535 5.565 125.905 6.065 ;
        RECT 126.185 5.565 126.555 6.065 ;
        RECT 127.485 5.565 127.855 6.065 ;
        RECT 128.135 5.565 128.505 6.065 ;
        RECT 129.435 5.565 129.805 6.065 ;
        RECT 130.085 5.565 130.455 6.065 ;
        RECT 131.385 5.565 131.755 6.065 ;
        RECT 132.035 5.565 132.405 6.065 ;
        RECT 133.335 5.565 133.705 6.065 ;
        RECT 133.985 5.565 134.355 6.065 ;
        RECT 135.285 5.565 135.655 6.065 ;
        RECT 64.115 3.585 65.115 3.985 ;
        RECT 68.235 3.585 69.235 3.985 ;
        RECT 72.135 3.585 73.135 3.985 ;
        RECT 76.035 3.585 77.035 3.985 ;
        RECT 122.075 3.585 123.075 3.985 ;
        RECT 126.195 3.585 127.195 3.985 ;
        RECT 130.095 3.585 131.095 3.985 ;
        RECT 133.995 3.585 134.995 3.985 ;
      LAYER met3 ;
        RECT 1.000 35.260 136.945 37.250 ;
        RECT 1.000 35.250 3.000 35.260 ;
        RECT 64.115 35.250 65.115 35.260 ;
        RECT 68.235 35.250 69.235 35.260 ;
        RECT 72.135 35.250 73.135 35.260 ;
        RECT 76.035 35.250 77.035 35.260 ;
        RECT 122.075 35.250 123.075 35.260 ;
        RECT 126.195 35.250 127.195 35.260 ;
        RECT 130.095 35.250 131.095 35.260 ;
        RECT 133.995 35.250 134.995 35.260 ;
        RECT 64.115 27.145 65.115 27.545 ;
        RECT 68.235 27.145 69.235 27.545 ;
        RECT 72.135 27.145 73.135 27.545 ;
        RECT 76.035 27.145 77.035 27.545 ;
        RECT 122.075 27.145 123.075 27.545 ;
        RECT 126.195 27.145 127.195 27.545 ;
        RECT 130.095 27.145 131.095 27.545 ;
        RECT 133.995 27.145 134.995 27.545 ;
        RECT 65.000 25.065 77.965 25.565 ;
        RECT 122.960 25.065 135.925 25.565 ;
        RECT 76.035 24.325 77.035 24.655 ;
        RECT 133.995 24.325 134.995 24.655 ;
        RECT 64.115 5.565 78.485 6.065 ;
        RECT 122.075 5.565 136.445 6.065 ;
        RECT 64.115 3.585 65.115 3.985 ;
        RECT 68.235 3.585 69.235 3.985 ;
        RECT 72.135 3.585 73.135 3.985 ;
        RECT 76.035 3.585 77.035 3.985 ;
        RECT 122.075 3.585 123.075 3.985 ;
        RECT 126.195 3.585 127.195 3.985 ;
        RECT 130.095 3.585 131.095 3.985 ;
        RECT 133.995 3.585 134.995 3.985 ;
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
        RECT 64.115 3.585 65.115 37.250 ;
        RECT 68.235 3.585 69.235 37.250 ;
        RECT 72.135 3.585 73.135 37.250 ;
        RECT 76.035 3.585 77.035 37.250 ;
        RECT 122.075 3.585 123.075 37.250 ;
        RECT 126.195 3.585 127.195 37.250 ;
        RECT 130.095 3.585 131.095 37.250 ;
        RECT 133.995 3.585 134.995 37.250 ;
    END
  END VDPWR
  PIN ua[1]
    ANTENNAGATEAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 122.940 16.065 123.270 16.395 ;
        RECT 124.580 16.145 124.910 16.315 ;
        RECT 126.530 16.145 126.860 16.315 ;
        RECT 128.480 16.145 128.810 16.315 ;
        RECT 130.430 16.145 130.760 16.315 ;
        RECT 132.380 16.145 132.710 16.315 ;
        RECT 124.580 14.815 124.910 14.985 ;
        RECT 126.530 14.815 126.860 14.985 ;
        RECT 128.480 14.815 128.810 14.985 ;
        RECT 130.430 14.815 130.760 14.985 ;
        RECT 132.380 14.815 132.710 14.985 ;
        RECT 134.330 14.815 134.660 14.985 ;
      LAYER met1 ;
        RECT 121.345 16.065 121.715 16.395 ;
        RECT 122.920 16.065 123.290 16.395 ;
        RECT 124.560 16.065 124.930 16.395 ;
        RECT 126.510 16.065 126.880 16.395 ;
        RECT 128.460 16.065 128.830 16.395 ;
        RECT 130.410 16.065 130.780 16.395 ;
        RECT 132.360 16.065 132.730 16.395 ;
        RECT 121.345 14.735 121.715 15.065 ;
        RECT 124.560 14.735 124.930 15.065 ;
        RECT 126.510 14.735 126.880 15.065 ;
        RECT 128.460 14.735 128.830 15.065 ;
        RECT 130.410 14.735 130.780 15.065 ;
        RECT 132.360 14.735 132.730 15.065 ;
        RECT 134.310 14.735 134.680 15.065 ;
      LAYER met2 ;
        RECT 121.345 16.065 121.715 16.395 ;
        RECT 122.920 16.065 123.290 16.395 ;
        RECT 124.560 16.065 124.930 16.395 ;
        RECT 126.510 16.065 126.880 16.395 ;
        RECT 128.460 16.065 128.830 16.395 ;
        RECT 130.410 16.065 130.780 16.395 ;
        RECT 132.360 16.065 132.730 16.395 ;
        RECT 121.395 15.065 121.665 16.065 ;
        RECT 121.345 14.735 121.715 15.065 ;
        RECT 124.560 14.735 124.930 15.065 ;
        RECT 126.510 14.735 126.880 15.065 ;
        RECT 128.460 14.735 128.830 15.065 ;
        RECT 130.410 14.735 130.780 15.065 ;
        RECT 132.360 14.735 132.730 15.065 ;
        RECT 134.310 14.735 134.680 15.065 ;
      LAYER met3 ;
        RECT 120.475 16.065 139.750 16.395 ;
        RECT 138.850 15.065 139.750 16.065 ;
        RECT 121.345 14.735 139.750 15.065 ;
      LAYER met4 ;
        RECT 138.850 2.400 139.750 16.395 ;
        RECT 132.490 1.500 139.750 2.400 ;
        RECT 132.490 0.000 133.390 1.500 ;
    END
  END ua[1]
  OBS
      LAYER li1 ;
        RECT 65.320 26.595 65.650 26.765 ;
        RECT 66.620 26.595 66.950 26.765 ;
        RECT 68.570 26.595 68.900 26.765 ;
        RECT 70.520 26.595 70.850 26.765 ;
        RECT 72.470 26.595 72.800 26.765 ;
        RECT 74.420 26.595 74.750 26.765 ;
        RECT 123.280 26.595 123.610 26.765 ;
        RECT 124.580 26.595 124.910 26.765 ;
        RECT 126.530 26.595 126.860 26.765 ;
        RECT 128.480 26.595 128.810 26.765 ;
        RECT 130.430 26.595 130.760 26.765 ;
        RECT 132.380 26.595 132.710 26.765 ;
        RECT 65.075 24.430 65.245 26.200 ;
        RECT 66.375 24.430 66.545 26.200 ;
        RECT 68.325 24.430 68.495 26.200 ;
        RECT 70.275 24.430 70.445 26.200 ;
        RECT 72.225 24.430 72.395 26.200 ;
        RECT 74.175 24.430 74.345 26.200 ;
        RECT 123.035 24.430 123.205 26.200 ;
        RECT 124.335 24.430 124.505 26.200 ;
        RECT 126.285 24.430 126.455 26.200 ;
        RECT 128.235 24.430 128.405 26.200 ;
        RECT 130.185 24.430 130.355 26.200 ;
        RECT 132.135 24.430 132.305 26.200 ;
        RECT 76.875 23.900 77.675 24.170 ;
        RECT 134.835 23.900 135.635 24.170 ;
        RECT 66.375 21.690 66.545 23.460 ;
        RECT 67.025 21.690 67.195 23.460 ;
        RECT 68.325 21.690 68.495 23.460 ;
        RECT 68.975 21.690 69.145 23.460 ;
        RECT 70.275 21.690 70.445 23.460 ;
        RECT 70.925 21.690 71.095 23.460 ;
        RECT 72.225 21.690 72.395 23.460 ;
        RECT 72.875 21.690 73.045 23.460 ;
        RECT 74.175 21.690 74.345 23.460 ;
        RECT 74.825 21.690 74.995 23.460 ;
        RECT 76.045 21.690 76.215 23.460 ;
        RECT 124.335 21.690 124.505 23.460 ;
        RECT 124.985 21.690 125.155 23.460 ;
        RECT 126.285 21.690 126.455 23.460 ;
        RECT 126.935 21.690 127.105 23.460 ;
        RECT 128.235 21.690 128.405 23.460 ;
        RECT 128.885 21.690 129.055 23.460 ;
        RECT 130.185 21.690 130.355 23.460 ;
        RECT 130.835 21.690 131.005 23.460 ;
        RECT 132.135 21.690 132.305 23.460 ;
        RECT 132.785 21.690 132.955 23.460 ;
        RECT 134.005 21.690 134.175 23.460 ;
        RECT 66.140 20.295 66.470 20.615 ;
        RECT 68.090 20.295 68.420 20.615 ;
        RECT 70.040 20.295 70.370 20.615 ;
        RECT 71.990 20.295 72.320 20.615 ;
        RECT 73.940 20.295 74.270 20.615 ;
        RECT 76.165 20.320 76.495 20.590 ;
        RECT 124.100 20.295 124.430 20.615 ;
        RECT 126.050 20.295 126.380 20.615 ;
        RECT 128.000 20.295 128.330 20.615 ;
        RECT 129.950 20.295 130.280 20.615 ;
        RECT 131.900 20.295 132.230 20.615 ;
        RECT 134.125 20.320 134.455 20.590 ;
        RECT 66.375 18.490 66.545 19.180 ;
        RECT 67.025 18.490 67.195 19.180 ;
        RECT 68.325 18.490 68.495 19.180 ;
        RECT 68.975 18.490 69.145 19.180 ;
        RECT 70.275 18.490 70.445 19.180 ;
        RECT 70.925 18.490 71.095 19.180 ;
        RECT 72.225 18.490 72.395 19.180 ;
        RECT 72.875 18.490 73.045 19.180 ;
        RECT 74.175 18.490 74.345 19.180 ;
        RECT 74.825 18.490 74.995 19.180 ;
        RECT 76.045 18.490 76.215 19.180 ;
        RECT 124.335 18.490 124.505 19.180 ;
        RECT 124.985 18.490 125.155 19.180 ;
        RECT 126.285 18.490 126.455 19.180 ;
        RECT 126.935 18.490 127.105 19.180 ;
        RECT 128.235 18.490 128.405 19.180 ;
        RECT 128.885 18.490 129.055 19.180 ;
        RECT 130.185 18.490 130.355 19.180 ;
        RECT 130.835 18.490 131.005 19.180 ;
        RECT 132.135 18.490 132.305 19.180 ;
        RECT 132.785 18.490 132.955 19.180 ;
        RECT 134.005 18.490 134.175 19.180 ;
        RECT 65.075 16.750 65.245 17.440 ;
        RECT 66.375 16.750 66.545 17.440 ;
        RECT 68.325 16.750 68.495 17.440 ;
        RECT 70.275 16.750 70.445 17.440 ;
        RECT 72.225 16.750 72.395 17.440 ;
        RECT 74.175 16.750 74.345 17.440 ;
        RECT 123.035 16.750 123.205 17.440 ;
        RECT 124.335 16.750 124.505 17.440 ;
        RECT 126.285 16.750 126.455 17.440 ;
        RECT 128.235 16.750 128.405 17.440 ;
        RECT 130.185 16.750 130.355 17.440 ;
        RECT 132.135 16.750 132.305 17.440 ;
        RECT 67.025 13.690 67.195 14.380 ;
        RECT 68.975 13.690 69.145 14.380 ;
        RECT 70.925 13.690 71.095 14.380 ;
        RECT 72.875 13.690 73.045 14.380 ;
        RECT 74.825 13.690 74.995 14.380 ;
        RECT 76.775 13.690 76.945 14.380 ;
        RECT 124.985 13.690 125.155 14.380 ;
        RECT 126.935 13.690 127.105 14.380 ;
        RECT 128.885 13.690 129.055 14.380 ;
        RECT 130.835 13.690 131.005 14.380 ;
        RECT 132.785 13.690 132.955 14.380 ;
        RECT 134.735 13.690 134.905 14.380 ;
        RECT 66.375 11.950 66.545 12.640 ;
        RECT 67.025 11.950 67.195 12.640 ;
        RECT 68.325 11.950 68.495 12.640 ;
        RECT 68.975 11.950 69.145 12.640 ;
        RECT 70.275 11.950 70.445 12.640 ;
        RECT 70.925 11.950 71.095 12.640 ;
        RECT 72.225 11.950 72.395 12.640 ;
        RECT 72.875 11.950 73.045 12.640 ;
        RECT 74.175 11.950 74.345 12.640 ;
        RECT 74.825 11.950 74.995 12.640 ;
        RECT 76.125 11.950 76.295 12.640 ;
        RECT 76.775 11.950 76.945 12.640 ;
        RECT 124.335 11.950 124.505 12.640 ;
        RECT 124.985 11.950 125.155 12.640 ;
        RECT 126.285 11.950 126.455 12.640 ;
        RECT 126.935 11.950 127.105 12.640 ;
        RECT 128.235 11.950 128.405 12.640 ;
        RECT 128.885 11.950 129.055 12.640 ;
        RECT 130.185 11.950 130.355 12.640 ;
        RECT 130.835 11.950 131.005 12.640 ;
        RECT 132.135 11.950 132.305 12.640 ;
        RECT 132.785 11.950 132.955 12.640 ;
        RECT 134.085 11.950 134.255 12.640 ;
        RECT 134.735 11.950 134.905 12.640 ;
        RECT 67.100 10.515 67.430 10.835 ;
        RECT 69.050 10.515 69.380 10.835 ;
        RECT 71.000 10.515 71.330 10.835 ;
        RECT 72.950 10.515 73.280 10.835 ;
        RECT 74.900 10.515 75.230 10.835 ;
        RECT 76.850 10.515 77.180 10.835 ;
        RECT 125.060 10.515 125.390 10.835 ;
        RECT 127.010 10.515 127.340 10.835 ;
        RECT 128.960 10.515 129.290 10.835 ;
        RECT 130.910 10.515 131.240 10.835 ;
        RECT 132.860 10.515 133.190 10.835 ;
        RECT 134.810 10.515 135.140 10.835 ;
        RECT 66.375 7.670 66.545 9.440 ;
        RECT 67.025 7.670 67.195 9.440 ;
        RECT 68.325 7.670 68.495 9.440 ;
        RECT 68.975 7.670 69.145 9.440 ;
        RECT 70.275 7.670 70.445 9.440 ;
        RECT 70.925 7.670 71.095 9.440 ;
        RECT 72.225 7.670 72.395 9.440 ;
        RECT 72.875 7.670 73.045 9.440 ;
        RECT 74.175 7.670 74.345 9.440 ;
        RECT 74.825 7.670 74.995 9.440 ;
        RECT 76.125 7.670 76.295 9.440 ;
        RECT 76.775 7.670 76.945 9.440 ;
        RECT 124.335 7.670 124.505 9.440 ;
        RECT 124.985 7.670 125.155 9.440 ;
        RECT 126.285 7.670 126.455 9.440 ;
        RECT 126.935 7.670 127.105 9.440 ;
        RECT 128.235 7.670 128.405 9.440 ;
        RECT 128.885 7.670 129.055 9.440 ;
        RECT 130.185 7.670 130.355 9.440 ;
        RECT 130.835 7.670 131.005 9.440 ;
        RECT 132.135 7.670 132.305 9.440 ;
        RECT 132.785 7.670 132.955 9.440 ;
        RECT 134.085 7.670 134.255 9.440 ;
        RECT 134.735 7.670 134.905 9.440 ;
        RECT 67.025 4.930 67.195 6.700 ;
        RECT 68.975 4.930 69.145 6.700 ;
        RECT 70.925 4.930 71.095 6.700 ;
        RECT 72.875 4.930 73.045 6.700 ;
        RECT 74.825 4.930 74.995 6.700 ;
        RECT 76.775 4.930 76.945 6.700 ;
        RECT 124.985 4.930 125.155 6.700 ;
        RECT 126.935 4.930 127.105 6.700 ;
        RECT 128.885 4.930 129.055 6.700 ;
        RECT 130.835 4.930 131.005 6.700 ;
        RECT 132.785 4.930 132.955 6.700 ;
        RECT 134.735 4.930 134.905 6.700 ;
        RECT 66.620 4.365 66.950 4.535 ;
        RECT 68.570 4.365 68.900 4.535 ;
        RECT 70.520 4.365 70.850 4.535 ;
        RECT 72.470 4.365 72.800 4.535 ;
        RECT 74.420 4.365 74.750 4.535 ;
        RECT 76.370 4.365 76.700 4.535 ;
        RECT 124.580 4.365 124.910 4.535 ;
        RECT 126.530 4.365 126.860 4.535 ;
        RECT 128.480 4.365 128.810 4.535 ;
        RECT 130.430 4.365 130.760 4.535 ;
        RECT 132.380 4.365 132.710 4.535 ;
        RECT 134.330 4.365 134.660 4.535 ;
      LAYER met1 ;
        RECT 62.465 26.515 62.835 26.845 ;
        RECT 65.000 26.515 65.670 26.845 ;
        RECT 66.600 26.515 66.970 26.845 ;
        RECT 68.550 26.515 68.920 26.845 ;
        RECT 70.500 26.515 70.870 26.845 ;
        RECT 72.450 26.515 72.820 26.845 ;
        RECT 74.400 26.515 74.770 26.845 ;
        RECT 120.425 26.515 120.795 26.845 ;
        RECT 122.960 26.515 123.630 26.845 ;
        RECT 124.560 26.515 124.930 26.845 ;
        RECT 126.510 26.515 126.880 26.845 ;
        RECT 128.460 26.515 128.830 26.845 ;
        RECT 130.410 26.515 130.780 26.845 ;
        RECT 132.360 26.515 132.730 26.845 ;
        RECT 65.000 24.450 65.320 26.180 ;
        RECT 66.345 21.710 66.575 26.180 ;
        RECT 66.950 21.710 67.270 23.440 ;
        RECT 68.295 21.710 68.525 26.180 ;
        RECT 68.900 21.710 69.220 23.440 ;
        RECT 70.245 21.710 70.475 26.180 ;
        RECT 70.850 21.710 71.170 23.440 ;
        RECT 72.195 21.710 72.425 26.180 ;
        RECT 72.800 21.710 73.120 23.440 ;
        RECT 74.145 21.710 74.375 26.180 ;
        RECT 122.960 24.450 123.280 26.180 ;
        RECT 75.990 24.135 76.310 24.165 ;
        RECT 76.875 24.135 77.675 24.170 ;
        RECT 75.990 23.935 77.675 24.135 ;
        RECT 75.990 23.905 76.310 23.935 ;
        RECT 76.875 23.900 77.675 23.935 ;
        RECT 74.750 21.710 75.070 23.440 ;
        RECT 76.015 21.985 76.245 23.440 ;
        RECT 75.970 21.725 76.290 21.985 ;
        RECT 76.015 21.710 76.245 21.725 ;
        RECT 124.305 21.710 124.535 26.180 ;
        RECT 124.910 21.710 125.230 23.440 ;
        RECT 126.255 21.710 126.485 26.180 ;
        RECT 126.860 21.710 127.180 23.440 ;
        RECT 128.205 21.710 128.435 26.180 ;
        RECT 128.810 21.710 129.130 23.440 ;
        RECT 130.155 21.710 130.385 26.180 ;
        RECT 130.760 21.710 131.080 23.440 ;
        RECT 132.105 21.710 132.335 26.180 ;
        RECT 133.950 24.135 134.270 24.165 ;
        RECT 134.835 24.135 135.635 24.170 ;
        RECT 133.950 23.935 135.635 24.135 ;
        RECT 133.950 23.905 134.270 23.935 ;
        RECT 134.835 23.900 135.635 23.935 ;
        RECT 132.710 21.710 133.030 23.440 ;
        RECT 133.975 21.985 134.205 23.440 ;
        RECT 133.930 21.725 134.250 21.985 ;
        RECT 133.975 21.710 134.205 21.725 ;
        RECT 64.455 20.295 66.470 20.615 ;
        RECT 66.950 20.295 68.420 20.615 ;
        RECT 68.900 20.295 70.370 20.615 ;
        RECT 70.850 20.295 72.320 20.615 ;
        RECT 72.800 20.295 74.270 20.615 ;
        RECT 74.750 20.295 78.645 20.615 ;
        RECT 122.415 20.295 124.430 20.615 ;
        RECT 124.910 20.295 126.380 20.615 ;
        RECT 126.860 20.295 128.330 20.615 ;
        RECT 128.810 20.295 130.280 20.615 ;
        RECT 130.760 20.295 132.230 20.615 ;
        RECT 132.710 20.295 136.605 20.615 ;
        RECT 65.000 16.770 65.320 17.420 ;
        RECT 66.345 16.770 66.575 19.160 ;
        RECT 66.950 18.510 67.270 19.160 ;
        RECT 68.295 16.770 68.525 19.160 ;
        RECT 68.900 18.510 69.220 19.160 ;
        RECT 70.245 16.770 70.475 19.160 ;
        RECT 70.850 18.510 71.170 19.160 ;
        RECT 72.195 16.770 72.425 19.160 ;
        RECT 72.800 18.510 73.120 19.160 ;
        RECT 74.145 16.770 74.375 19.160 ;
        RECT 74.750 18.510 75.070 19.160 ;
        RECT 76.015 19.145 76.245 19.160 ;
        RECT 75.970 18.885 76.290 19.145 ;
        RECT 76.015 18.510 76.245 18.885 ;
        RECT 122.960 16.770 123.280 17.420 ;
        RECT 124.305 16.770 124.535 19.160 ;
        RECT 124.910 18.510 125.230 19.160 ;
        RECT 126.255 16.770 126.485 19.160 ;
        RECT 126.860 18.510 127.180 19.160 ;
        RECT 128.205 16.770 128.435 19.160 ;
        RECT 128.810 18.510 129.130 19.160 ;
        RECT 130.155 16.770 130.385 19.160 ;
        RECT 130.760 18.510 131.080 19.160 ;
        RECT 132.105 16.770 132.335 19.160 ;
        RECT 132.710 18.510 133.030 19.160 ;
        RECT 133.975 19.145 134.205 19.160 ;
        RECT 133.930 18.885 134.250 19.145 ;
        RECT 133.975 18.510 134.205 18.885 ;
        RECT 66.300 11.970 66.620 12.620 ;
        RECT 66.995 11.970 67.225 14.360 ;
        RECT 68.250 11.970 68.570 12.620 ;
        RECT 68.945 11.970 69.175 14.360 ;
        RECT 70.200 11.970 70.520 12.620 ;
        RECT 70.895 11.970 71.125 14.360 ;
        RECT 72.150 11.970 72.470 12.620 ;
        RECT 72.845 11.970 73.075 14.360 ;
        RECT 74.100 11.970 74.420 12.620 ;
        RECT 74.795 11.970 75.025 14.360 ;
        RECT 76.050 11.970 76.370 12.620 ;
        RECT 76.745 11.970 76.975 14.360 ;
        RECT 124.260 11.970 124.580 12.620 ;
        RECT 124.955 11.970 125.185 14.360 ;
        RECT 126.210 11.970 126.530 12.620 ;
        RECT 126.905 11.970 127.135 14.360 ;
        RECT 128.160 11.970 128.480 12.620 ;
        RECT 128.855 11.970 129.085 14.360 ;
        RECT 130.110 11.970 130.430 12.620 ;
        RECT 130.805 11.970 131.035 14.360 ;
        RECT 132.060 11.970 132.380 12.620 ;
        RECT 132.755 11.970 132.985 14.360 ;
        RECT 134.010 11.970 134.330 12.620 ;
        RECT 134.705 11.970 134.935 14.360 ;
        RECT 64.455 10.515 66.620 10.835 ;
        RECT 67.100 10.515 68.570 10.835 ;
        RECT 69.050 10.515 70.520 10.835 ;
        RECT 71.000 10.515 72.470 10.835 ;
        RECT 72.950 10.515 74.420 10.835 ;
        RECT 74.900 10.515 76.370 10.835 ;
        RECT 76.850 10.515 78.645 10.835 ;
        RECT 122.415 10.515 124.580 10.835 ;
        RECT 125.060 10.515 126.530 10.835 ;
        RECT 127.010 10.515 128.480 10.835 ;
        RECT 128.960 10.515 130.430 10.835 ;
        RECT 130.910 10.515 132.380 10.835 ;
        RECT 132.860 10.515 134.330 10.835 ;
        RECT 134.810 10.515 136.605 10.835 ;
        RECT 66.300 7.690 66.620 9.420 ;
        RECT 66.995 4.950 67.225 9.420 ;
        RECT 68.250 7.690 68.570 9.420 ;
        RECT 68.945 4.950 69.175 9.420 ;
        RECT 70.200 7.690 70.520 9.420 ;
        RECT 70.895 4.950 71.125 9.420 ;
        RECT 72.150 7.690 72.470 9.420 ;
        RECT 72.845 4.950 73.075 9.420 ;
        RECT 74.100 7.690 74.420 9.420 ;
        RECT 74.795 4.950 75.025 9.420 ;
        RECT 76.050 7.690 76.370 9.420 ;
        RECT 76.745 4.950 76.975 9.420 ;
        RECT 124.260 7.690 124.580 9.420 ;
        RECT 124.955 4.950 125.185 9.420 ;
        RECT 126.210 7.690 126.530 9.420 ;
        RECT 126.905 4.950 127.135 9.420 ;
        RECT 128.160 7.690 128.480 9.420 ;
        RECT 128.855 4.950 129.085 9.420 ;
        RECT 130.110 7.690 130.430 9.420 ;
        RECT 130.805 4.950 131.035 9.420 ;
        RECT 132.060 7.690 132.380 9.420 ;
        RECT 132.755 4.950 132.985 9.420 ;
        RECT 134.010 7.690 134.330 9.420 ;
        RECT 134.705 4.950 134.935 9.420 ;
        RECT 62.465 4.285 62.835 4.615 ;
        RECT 66.600 4.285 66.970 4.615 ;
        RECT 68.550 4.285 68.920 4.615 ;
        RECT 70.500 4.285 70.870 4.615 ;
        RECT 72.450 4.285 72.820 4.615 ;
        RECT 74.400 4.285 74.770 4.615 ;
        RECT 76.350 4.285 76.720 4.615 ;
        RECT 120.425 4.285 120.795 4.615 ;
        RECT 124.560 4.285 124.930 4.615 ;
        RECT 126.510 4.285 126.880 4.615 ;
        RECT 128.460 4.285 128.830 4.615 ;
        RECT 130.410 4.285 130.780 4.615 ;
        RECT 132.360 4.285 132.730 4.615 ;
        RECT 134.310 4.285 134.680 4.615 ;
      LAYER met2 ;
        RECT 62.465 26.515 62.835 26.845 ;
        RECT 65.000 26.515 65.670 26.845 ;
        RECT 66.600 26.515 66.970 26.845 ;
        RECT 68.550 26.515 68.920 26.845 ;
        RECT 70.500 26.515 70.870 26.845 ;
        RECT 72.450 26.515 72.820 26.845 ;
        RECT 74.400 26.515 74.770 26.845 ;
        RECT 120.425 26.515 120.795 26.845 ;
        RECT 122.960 26.515 123.630 26.845 ;
        RECT 124.560 26.515 124.930 26.845 ;
        RECT 126.510 26.515 126.880 26.845 ;
        RECT 128.460 26.515 128.830 26.845 ;
        RECT 130.410 26.515 130.780 26.845 ;
        RECT 132.360 26.515 132.730 26.845 ;
        RECT 62.515 4.615 62.785 26.515 ;
        RECT 64.455 10.515 64.775 20.615 ;
        RECT 65.000 16.770 65.320 26.515 ;
        RECT 75.990 23.905 76.310 24.165 ;
        RECT 66.950 21.710 67.270 23.440 ;
        RECT 68.900 21.710 69.220 23.440 ;
        RECT 70.850 21.710 71.170 23.440 ;
        RECT 72.800 21.710 73.120 23.440 ;
        RECT 74.750 21.710 75.070 23.440 ;
        RECT 76.025 21.985 76.225 23.905 ;
        RECT 75.970 21.725 76.290 21.985 ;
        RECT 66.995 20.615 67.225 21.710 ;
        RECT 68.945 20.615 69.175 21.710 ;
        RECT 70.895 20.615 71.125 21.710 ;
        RECT 72.845 20.615 73.075 21.710 ;
        RECT 74.795 20.615 75.025 21.710 ;
        RECT 66.950 20.295 67.270 20.615 ;
        RECT 68.900 20.295 69.220 20.615 ;
        RECT 70.850 20.295 71.170 20.615 ;
        RECT 72.800 20.295 73.120 20.615 ;
        RECT 74.750 20.295 75.070 20.615 ;
        RECT 66.995 19.160 67.225 20.295 ;
        RECT 68.945 19.160 69.175 20.295 ;
        RECT 70.895 19.160 71.125 20.295 ;
        RECT 72.845 19.160 73.075 20.295 ;
        RECT 74.795 19.160 75.025 20.295 ;
        RECT 66.950 18.510 67.270 19.160 ;
        RECT 68.900 18.510 69.220 19.160 ;
        RECT 70.850 18.510 71.170 19.160 ;
        RECT 72.800 18.510 73.120 19.160 ;
        RECT 74.750 18.510 75.070 19.160 ;
        RECT 76.025 19.145 76.225 21.725 ;
        RECT 75.970 18.885 76.290 19.145 ;
        RECT 66.300 11.970 66.620 12.620 ;
        RECT 68.250 11.970 68.570 12.620 ;
        RECT 70.200 11.970 70.520 12.620 ;
        RECT 72.150 11.970 72.470 12.620 ;
        RECT 74.100 11.970 74.420 12.620 ;
        RECT 76.050 11.970 76.370 12.620 ;
        RECT 66.345 10.835 66.575 11.970 ;
        RECT 68.295 10.835 68.525 11.970 ;
        RECT 70.245 10.835 70.475 11.970 ;
        RECT 72.195 10.835 72.425 11.970 ;
        RECT 74.145 10.835 74.375 11.970 ;
        RECT 76.095 10.835 76.325 11.970 ;
        RECT 66.300 10.515 66.620 10.835 ;
        RECT 68.250 10.515 68.570 10.835 ;
        RECT 70.200 10.515 70.520 10.835 ;
        RECT 72.150 10.515 72.470 10.835 ;
        RECT 74.100 10.515 74.420 10.835 ;
        RECT 76.050 10.515 76.370 10.835 ;
        RECT 78.325 10.515 78.645 20.615 ;
        RECT 66.345 9.420 66.575 10.515 ;
        RECT 68.295 9.420 68.525 10.515 ;
        RECT 70.245 9.420 70.475 10.515 ;
        RECT 72.195 9.420 72.425 10.515 ;
        RECT 74.145 9.420 74.375 10.515 ;
        RECT 76.095 9.420 76.325 10.515 ;
        RECT 66.300 7.690 66.620 9.420 ;
        RECT 68.250 7.690 68.570 9.420 ;
        RECT 70.200 7.690 70.520 9.420 ;
        RECT 72.150 7.690 72.470 9.420 ;
        RECT 74.100 7.690 74.420 9.420 ;
        RECT 76.050 7.690 76.370 9.420 ;
        RECT 120.475 4.615 120.745 26.515 ;
        RECT 122.415 10.515 122.735 20.615 ;
        RECT 122.960 16.770 123.280 26.515 ;
        RECT 133.950 23.905 134.270 24.165 ;
        RECT 124.910 21.710 125.230 23.440 ;
        RECT 126.860 21.710 127.180 23.440 ;
        RECT 128.810 21.710 129.130 23.440 ;
        RECT 130.760 21.710 131.080 23.440 ;
        RECT 132.710 21.710 133.030 23.440 ;
        RECT 133.985 21.985 134.185 23.905 ;
        RECT 133.930 21.725 134.250 21.985 ;
        RECT 124.955 20.615 125.185 21.710 ;
        RECT 126.905 20.615 127.135 21.710 ;
        RECT 128.855 20.615 129.085 21.710 ;
        RECT 130.805 20.615 131.035 21.710 ;
        RECT 132.755 20.615 132.985 21.710 ;
        RECT 124.910 20.295 125.230 20.615 ;
        RECT 126.860 20.295 127.180 20.615 ;
        RECT 128.810 20.295 129.130 20.615 ;
        RECT 130.760 20.295 131.080 20.615 ;
        RECT 132.710 20.295 133.030 20.615 ;
        RECT 124.955 19.160 125.185 20.295 ;
        RECT 126.905 19.160 127.135 20.295 ;
        RECT 128.855 19.160 129.085 20.295 ;
        RECT 130.805 19.160 131.035 20.295 ;
        RECT 132.755 19.160 132.985 20.295 ;
        RECT 124.910 18.510 125.230 19.160 ;
        RECT 126.860 18.510 127.180 19.160 ;
        RECT 128.810 18.510 129.130 19.160 ;
        RECT 130.760 18.510 131.080 19.160 ;
        RECT 132.710 18.510 133.030 19.160 ;
        RECT 133.985 19.145 134.185 21.725 ;
        RECT 133.930 18.885 134.250 19.145 ;
        RECT 124.260 11.970 124.580 12.620 ;
        RECT 126.210 11.970 126.530 12.620 ;
        RECT 128.160 11.970 128.480 12.620 ;
        RECT 130.110 11.970 130.430 12.620 ;
        RECT 132.060 11.970 132.380 12.620 ;
        RECT 134.010 11.970 134.330 12.620 ;
        RECT 124.305 10.835 124.535 11.970 ;
        RECT 126.255 10.835 126.485 11.970 ;
        RECT 128.205 10.835 128.435 11.970 ;
        RECT 130.155 10.835 130.385 11.970 ;
        RECT 132.105 10.835 132.335 11.970 ;
        RECT 134.055 10.835 134.285 11.970 ;
        RECT 124.260 10.515 124.580 10.835 ;
        RECT 126.210 10.515 126.530 10.835 ;
        RECT 128.160 10.515 128.480 10.835 ;
        RECT 130.110 10.515 130.430 10.835 ;
        RECT 132.060 10.515 132.380 10.835 ;
        RECT 134.010 10.515 134.330 10.835 ;
        RECT 136.285 10.515 136.605 20.615 ;
        RECT 124.305 9.420 124.535 10.515 ;
        RECT 126.255 9.420 126.485 10.515 ;
        RECT 128.205 9.420 128.435 10.515 ;
        RECT 130.155 9.420 130.385 10.515 ;
        RECT 132.105 9.420 132.335 10.515 ;
        RECT 134.055 9.420 134.285 10.515 ;
        RECT 124.260 7.690 124.580 9.420 ;
        RECT 126.210 7.690 126.530 9.420 ;
        RECT 128.160 7.690 128.480 9.420 ;
        RECT 130.110 7.690 130.430 9.420 ;
        RECT 132.060 7.690 132.380 9.420 ;
        RECT 134.010 7.690 134.330 9.420 ;
        RECT 62.465 4.285 62.835 4.615 ;
        RECT 66.600 4.285 66.970 4.615 ;
        RECT 68.550 4.285 68.920 4.615 ;
        RECT 70.500 4.285 70.870 4.615 ;
        RECT 72.450 4.285 72.820 4.615 ;
        RECT 74.400 4.285 74.770 4.615 ;
        RECT 76.350 4.285 76.720 4.615 ;
        RECT 120.425 4.285 120.795 4.615 ;
        RECT 124.560 4.285 124.930 4.615 ;
        RECT 126.510 4.285 126.880 4.615 ;
        RECT 128.460 4.285 128.830 4.615 ;
        RECT 130.410 4.285 130.780 4.615 ;
        RECT 132.360 4.285 132.730 4.615 ;
        RECT 134.310 4.285 134.680 4.615 ;
      LAYER met3 ;
        RECT 62.465 26.515 77.965 26.845 ;
        RECT 120.425 26.515 135.925 26.845 ;
        RECT 62.465 4.285 78.485 4.615 ;
        RECT 120.425 4.285 136.445 4.615 ;
  END
END tt_um_Onchip_VCOx2
END LIBRARY

