magic
tech sky130A
magscale 1 2
timestamp 1762792651
<< nwell >>
rect 12941 4791 15593 5545
rect 24533 4791 27185 5545
rect 12941 4239 15677 4791
rect 24533 4239 27269 4791
rect 12941 4171 15593 4239
rect 24533 4171 27185 4239
rect 12941 681 15593 2055
rect 24533 681 27185 2055
<< pwell >>
rect 13236 3641 15642 3893
rect 24828 3641 27234 3893
rect 13236 3545 15553 3641
rect 24828 3545 27145 3641
rect 12976 3507 15553 3545
rect 24568 3507 27145 3545
rect 12976 3179 15168 3507
rect 24568 3179 26760 3507
rect 12972 3047 15528 3179
rect 24564 3047 27120 3179
rect 13106 2933 15528 3047
rect 24698 2933 27120 3047
rect 13106 2681 15558 2933
rect 24698 2681 27150 2933
rect 13106 2333 15428 2681
rect 24698 2333 27020 2681
<< nmos >>
rect 15256 3667 15286 3867
rect 15346 3667 15376 3867
rect 15436 3667 15466 3867
rect 15526 3667 15556 3867
rect 26848 3667 26878 3867
rect 26938 3667 26968 3867
rect 27028 3667 27058 3867
rect 27118 3667 27148 3867
<< pmos >>
rect 15256 4315 15286 4715
rect 15346 4315 15376 4715
rect 15436 4315 15466 4715
rect 15526 4315 15556 4715
rect 26848 4315 26878 4715
rect 26938 4315 26968 4715
rect 27028 4315 27058 4715
rect 27118 4315 27148 4715
<< pmoslvt >>
rect 13062 4863 13132 5263
rect 13192 4863 13262 5263
rect 13322 4863 13392 5263
rect 13452 4863 13522 5263
rect 13582 4863 13652 5263
rect 13712 4863 13782 5263
rect 13842 4863 13912 5263
rect 13972 4863 14042 5263
rect 14102 4863 14172 5263
rect 14232 4863 14302 5263
rect 14362 4863 14432 5263
rect 14492 4863 14562 5263
rect 14622 4863 14692 5263
rect 14752 4863 14822 5263
rect 14882 4863 14952 5263
rect 15012 4863 15082 5263
rect 24654 4863 24724 5263
rect 24784 4863 24854 5263
rect 24914 4863 24984 5263
rect 25044 4863 25114 5263
rect 25174 4863 25244 5263
rect 25304 4863 25374 5263
rect 25434 4863 25504 5263
rect 25564 4863 25634 5263
rect 25694 4863 25764 5263
rect 25824 4863 25894 5263
rect 25954 4863 26024 5263
rect 26084 4863 26154 5263
rect 26214 4863 26284 5263
rect 26344 4863 26414 5263
rect 26474 4863 26544 5263
rect 26604 4863 26674 5263
rect 13322 4315 13392 4715
rect 13712 4315 13782 4715
rect 14102 4315 14172 4715
rect 14492 4315 14562 4715
rect 14882 4315 14952 4715
rect 24914 4315 24984 4715
rect 25304 4315 25374 4715
rect 25694 4315 25764 4715
rect 26084 4315 26154 4715
rect 26474 4315 26544 4715
rect 13322 1511 13392 1911
rect 13712 1511 13782 1911
rect 14102 1511 14172 1911
rect 14492 1511 14562 1911
rect 14882 1511 14952 1911
rect 15272 1511 15342 1911
rect 24914 1511 24984 1911
rect 25304 1511 25374 1911
rect 25694 1511 25764 1911
rect 26084 1511 26154 1911
rect 26474 1511 26544 1911
rect 26864 1511 26934 1911
rect 13192 963 13262 1363
rect 13322 963 13392 1363
rect 13452 963 13522 1363
rect 13582 963 13652 1363
rect 13712 963 13782 1363
rect 13842 963 13912 1363
rect 13972 963 14042 1363
rect 14102 963 14172 1363
rect 14232 963 14302 1363
rect 14362 963 14432 1363
rect 14492 963 14562 1363
rect 14622 963 14692 1363
rect 14752 963 14822 1363
rect 14882 963 14952 1363
rect 15012 963 15082 1363
rect 15142 963 15212 1363
rect 15272 963 15342 1363
rect 15402 963 15472 1363
rect 24784 963 24854 1363
rect 24914 963 24984 1363
rect 25044 963 25114 1363
rect 25174 963 25244 1363
rect 25304 963 25374 1363
rect 25434 963 25504 1363
rect 25564 963 25634 1363
rect 25694 963 25764 1363
rect 25824 963 25894 1363
rect 25954 963 26024 1363
rect 26084 963 26154 1363
rect 26214 963 26284 1363
rect 26344 963 26414 1363
rect 26474 963 26544 1363
rect 26604 963 26674 1363
rect 26734 963 26804 1363
rect 26864 963 26934 1363
rect 26994 963 27064 1363
<< nmoslvt >>
rect 13322 3667 13392 3867
rect 13452 3667 13522 3867
rect 13712 3667 13782 3867
rect 13842 3667 13912 3867
rect 14102 3667 14172 3867
rect 14232 3667 14302 3867
rect 14492 3667 14562 3867
rect 14622 3667 14692 3867
rect 14882 3667 14952 3867
rect 15012 3667 15082 3867
rect 24914 3667 24984 3867
rect 25044 3667 25114 3867
rect 25304 3667 25374 3867
rect 25434 3667 25504 3867
rect 25694 3667 25764 3867
rect 25824 3667 25894 3867
rect 26084 3667 26154 3867
rect 26214 3667 26284 3867
rect 26474 3667 26544 3867
rect 26604 3667 26674 3867
rect 13062 3319 13132 3519
rect 13192 3319 13262 3519
rect 13322 3319 13392 3519
rect 13452 3319 13522 3519
rect 13582 3319 13652 3519
rect 13712 3319 13782 3519
rect 13842 3319 13912 3519
rect 13972 3319 14042 3519
rect 14102 3319 14172 3519
rect 14232 3319 14302 3519
rect 14362 3319 14432 3519
rect 14492 3319 14562 3519
rect 14622 3319 14692 3519
rect 14752 3319 14822 3519
rect 14882 3319 14952 3519
rect 15012 3319 15082 3519
rect 24654 3319 24724 3519
rect 24784 3319 24854 3519
rect 24914 3319 24984 3519
rect 25044 3319 25114 3519
rect 25174 3319 25244 3519
rect 25304 3319 25374 3519
rect 25434 3319 25504 3519
rect 25564 3319 25634 3519
rect 25694 3319 25764 3519
rect 25824 3319 25894 3519
rect 25954 3319 26024 3519
rect 26084 3319 26154 3519
rect 26214 3319 26284 3519
rect 26344 3319 26414 3519
rect 26474 3319 26544 3519
rect 26604 3319 26674 3519
rect 13192 2707 13262 2907
rect 13322 2707 13392 2907
rect 13452 2707 13522 2907
rect 13582 2707 13652 2907
rect 13712 2707 13782 2907
rect 13842 2707 13912 2907
rect 13972 2707 14042 2907
rect 14102 2707 14172 2907
rect 14232 2707 14302 2907
rect 14362 2707 14432 2907
rect 14492 2707 14562 2907
rect 14622 2707 14692 2907
rect 14752 2707 14822 2907
rect 14882 2707 14952 2907
rect 15012 2707 15082 2907
rect 15142 2707 15212 2907
rect 15272 2707 15342 2907
rect 15402 2707 15472 2907
rect 24784 2707 24854 2907
rect 24914 2707 24984 2907
rect 25044 2707 25114 2907
rect 25174 2707 25244 2907
rect 25304 2707 25374 2907
rect 25434 2707 25504 2907
rect 25564 2707 25634 2907
rect 25694 2707 25764 2907
rect 25824 2707 25894 2907
rect 25954 2707 26024 2907
rect 26084 2707 26154 2907
rect 26214 2707 26284 2907
rect 26344 2707 26414 2907
rect 26474 2707 26544 2907
rect 26604 2707 26674 2907
rect 26734 2707 26804 2907
rect 26864 2707 26934 2907
rect 26994 2707 27064 2907
rect 13192 2359 13262 2559
rect 13322 2359 13392 2559
rect 13582 2359 13652 2559
rect 13712 2359 13782 2559
rect 13972 2359 14042 2559
rect 14102 2359 14172 2559
rect 14362 2359 14432 2559
rect 14492 2359 14562 2559
rect 14752 2359 14822 2559
rect 14882 2359 14952 2559
rect 15142 2359 15212 2559
rect 15272 2359 15342 2559
rect 24784 2359 24854 2559
rect 24914 2359 24984 2559
rect 25174 2359 25244 2559
rect 25304 2359 25374 2559
rect 25564 2359 25634 2559
rect 25694 2359 25764 2559
rect 25954 2359 26024 2559
rect 26084 2359 26154 2559
rect 26344 2359 26414 2559
rect 26474 2359 26544 2559
rect 26734 2359 26804 2559
rect 26864 2359 26934 2559
<< ndiff >>
rect 13262 3820 13322 3867
rect 13262 3786 13275 3820
rect 13309 3786 13322 3820
rect 13262 3748 13322 3786
rect 13262 3714 13275 3748
rect 13309 3714 13322 3748
rect 13262 3667 13322 3714
rect 13392 3820 13452 3867
rect 13392 3786 13405 3820
rect 13439 3786 13452 3820
rect 13392 3748 13452 3786
rect 13392 3714 13405 3748
rect 13439 3714 13452 3748
rect 13392 3667 13452 3714
rect 13522 3820 13582 3867
rect 13522 3786 13535 3820
rect 13569 3786 13582 3820
rect 13522 3748 13582 3786
rect 13522 3714 13535 3748
rect 13569 3714 13582 3748
rect 13522 3667 13582 3714
rect 13652 3820 13712 3867
rect 13652 3786 13665 3820
rect 13699 3786 13712 3820
rect 13652 3748 13712 3786
rect 13652 3714 13665 3748
rect 13699 3714 13712 3748
rect 13652 3667 13712 3714
rect 13782 3820 13842 3867
rect 13782 3786 13795 3820
rect 13829 3786 13842 3820
rect 13782 3748 13842 3786
rect 13782 3714 13795 3748
rect 13829 3714 13842 3748
rect 13782 3667 13842 3714
rect 13912 3820 13972 3867
rect 13912 3786 13925 3820
rect 13959 3786 13972 3820
rect 13912 3748 13972 3786
rect 13912 3714 13925 3748
rect 13959 3714 13972 3748
rect 13912 3667 13972 3714
rect 14042 3820 14102 3867
rect 14042 3786 14055 3820
rect 14089 3786 14102 3820
rect 14042 3748 14102 3786
rect 14042 3714 14055 3748
rect 14089 3714 14102 3748
rect 14042 3667 14102 3714
rect 14172 3820 14232 3867
rect 14172 3786 14185 3820
rect 14219 3786 14232 3820
rect 14172 3748 14232 3786
rect 14172 3714 14185 3748
rect 14219 3714 14232 3748
rect 14172 3667 14232 3714
rect 14302 3820 14362 3867
rect 14302 3786 14315 3820
rect 14349 3786 14362 3820
rect 14302 3748 14362 3786
rect 14302 3714 14315 3748
rect 14349 3714 14362 3748
rect 14302 3667 14362 3714
rect 14432 3820 14492 3867
rect 14432 3786 14445 3820
rect 14479 3786 14492 3820
rect 14432 3748 14492 3786
rect 14432 3714 14445 3748
rect 14479 3714 14492 3748
rect 14432 3667 14492 3714
rect 14562 3820 14622 3867
rect 14562 3786 14575 3820
rect 14609 3786 14622 3820
rect 14562 3748 14622 3786
rect 14562 3714 14575 3748
rect 14609 3714 14622 3748
rect 14562 3667 14622 3714
rect 14692 3820 14752 3867
rect 14692 3786 14705 3820
rect 14739 3786 14752 3820
rect 14692 3748 14752 3786
rect 14692 3714 14705 3748
rect 14739 3714 14752 3748
rect 14692 3667 14752 3714
rect 14822 3820 14882 3867
rect 14822 3786 14835 3820
rect 14869 3786 14882 3820
rect 14822 3748 14882 3786
rect 14822 3714 14835 3748
rect 14869 3714 14882 3748
rect 14822 3667 14882 3714
rect 14952 3820 15012 3867
rect 14952 3786 14965 3820
rect 14999 3786 15012 3820
rect 14952 3748 15012 3786
rect 14952 3714 14965 3748
rect 14999 3714 15012 3748
rect 14952 3667 15012 3714
rect 15082 3820 15142 3867
rect 15082 3786 15095 3820
rect 15129 3786 15142 3820
rect 15082 3748 15142 3786
rect 15082 3714 15095 3748
rect 15129 3714 15142 3748
rect 15082 3667 15142 3714
rect 15196 3820 15256 3867
rect 15196 3786 15209 3820
rect 15243 3786 15256 3820
rect 15196 3748 15256 3786
rect 15196 3714 15209 3748
rect 15243 3714 15256 3748
rect 15196 3667 15256 3714
rect 15286 3820 15346 3867
rect 15286 3786 15299 3820
rect 15333 3786 15346 3820
rect 15286 3748 15346 3786
rect 15286 3714 15299 3748
rect 15333 3714 15346 3748
rect 15286 3667 15346 3714
rect 15376 3820 15436 3867
rect 15376 3786 15389 3820
rect 15423 3786 15436 3820
rect 15376 3748 15436 3786
rect 15376 3714 15389 3748
rect 15423 3714 15436 3748
rect 15376 3667 15436 3714
rect 15466 3820 15526 3867
rect 15466 3786 15479 3820
rect 15513 3786 15526 3820
rect 15466 3748 15526 3786
rect 15466 3714 15479 3748
rect 15513 3714 15526 3748
rect 15466 3667 15526 3714
rect 15556 3820 15616 3867
rect 15556 3786 15569 3820
rect 15603 3786 15616 3820
rect 15556 3748 15616 3786
rect 15556 3714 15569 3748
rect 15603 3714 15616 3748
rect 15556 3667 15616 3714
rect 24854 3820 24914 3867
rect 24854 3786 24867 3820
rect 24901 3786 24914 3820
rect 24854 3748 24914 3786
rect 24854 3714 24867 3748
rect 24901 3714 24914 3748
rect 24854 3667 24914 3714
rect 24984 3820 25044 3867
rect 24984 3786 24997 3820
rect 25031 3786 25044 3820
rect 24984 3748 25044 3786
rect 24984 3714 24997 3748
rect 25031 3714 25044 3748
rect 24984 3667 25044 3714
rect 25114 3820 25174 3867
rect 25114 3786 25127 3820
rect 25161 3786 25174 3820
rect 25114 3748 25174 3786
rect 25114 3714 25127 3748
rect 25161 3714 25174 3748
rect 25114 3667 25174 3714
rect 25244 3820 25304 3867
rect 25244 3786 25257 3820
rect 25291 3786 25304 3820
rect 25244 3748 25304 3786
rect 25244 3714 25257 3748
rect 25291 3714 25304 3748
rect 25244 3667 25304 3714
rect 25374 3820 25434 3867
rect 25374 3786 25387 3820
rect 25421 3786 25434 3820
rect 25374 3748 25434 3786
rect 25374 3714 25387 3748
rect 25421 3714 25434 3748
rect 25374 3667 25434 3714
rect 25504 3820 25564 3867
rect 25504 3786 25517 3820
rect 25551 3786 25564 3820
rect 25504 3748 25564 3786
rect 25504 3714 25517 3748
rect 25551 3714 25564 3748
rect 25504 3667 25564 3714
rect 25634 3820 25694 3867
rect 25634 3786 25647 3820
rect 25681 3786 25694 3820
rect 25634 3748 25694 3786
rect 25634 3714 25647 3748
rect 25681 3714 25694 3748
rect 25634 3667 25694 3714
rect 25764 3820 25824 3867
rect 25764 3786 25777 3820
rect 25811 3786 25824 3820
rect 25764 3748 25824 3786
rect 25764 3714 25777 3748
rect 25811 3714 25824 3748
rect 25764 3667 25824 3714
rect 25894 3820 25954 3867
rect 25894 3786 25907 3820
rect 25941 3786 25954 3820
rect 25894 3748 25954 3786
rect 25894 3714 25907 3748
rect 25941 3714 25954 3748
rect 25894 3667 25954 3714
rect 26024 3820 26084 3867
rect 26024 3786 26037 3820
rect 26071 3786 26084 3820
rect 26024 3748 26084 3786
rect 26024 3714 26037 3748
rect 26071 3714 26084 3748
rect 26024 3667 26084 3714
rect 26154 3820 26214 3867
rect 26154 3786 26167 3820
rect 26201 3786 26214 3820
rect 26154 3748 26214 3786
rect 26154 3714 26167 3748
rect 26201 3714 26214 3748
rect 26154 3667 26214 3714
rect 26284 3820 26344 3867
rect 26284 3786 26297 3820
rect 26331 3786 26344 3820
rect 26284 3748 26344 3786
rect 26284 3714 26297 3748
rect 26331 3714 26344 3748
rect 26284 3667 26344 3714
rect 26414 3820 26474 3867
rect 26414 3786 26427 3820
rect 26461 3786 26474 3820
rect 26414 3748 26474 3786
rect 26414 3714 26427 3748
rect 26461 3714 26474 3748
rect 26414 3667 26474 3714
rect 26544 3820 26604 3867
rect 26544 3786 26557 3820
rect 26591 3786 26604 3820
rect 26544 3748 26604 3786
rect 26544 3714 26557 3748
rect 26591 3714 26604 3748
rect 26544 3667 26604 3714
rect 26674 3820 26734 3867
rect 26674 3786 26687 3820
rect 26721 3786 26734 3820
rect 26674 3748 26734 3786
rect 26674 3714 26687 3748
rect 26721 3714 26734 3748
rect 26674 3667 26734 3714
rect 26788 3820 26848 3867
rect 26788 3786 26801 3820
rect 26835 3786 26848 3820
rect 26788 3748 26848 3786
rect 26788 3714 26801 3748
rect 26835 3714 26848 3748
rect 26788 3667 26848 3714
rect 26878 3820 26938 3867
rect 26878 3786 26891 3820
rect 26925 3786 26938 3820
rect 26878 3748 26938 3786
rect 26878 3714 26891 3748
rect 26925 3714 26938 3748
rect 26878 3667 26938 3714
rect 26968 3820 27028 3867
rect 26968 3786 26981 3820
rect 27015 3786 27028 3820
rect 26968 3748 27028 3786
rect 26968 3714 26981 3748
rect 27015 3714 27028 3748
rect 26968 3667 27028 3714
rect 27058 3820 27118 3867
rect 27058 3786 27071 3820
rect 27105 3786 27118 3820
rect 27058 3748 27118 3786
rect 27058 3714 27071 3748
rect 27105 3714 27118 3748
rect 27058 3667 27118 3714
rect 27148 3820 27208 3867
rect 27148 3786 27161 3820
rect 27195 3786 27208 3820
rect 27148 3748 27208 3786
rect 27148 3714 27161 3748
rect 27195 3714 27208 3748
rect 27148 3667 27208 3714
rect 13002 3472 13062 3519
rect 13002 3438 13015 3472
rect 13049 3438 13062 3472
rect 13002 3400 13062 3438
rect 13002 3366 13015 3400
rect 13049 3366 13062 3400
rect 13002 3319 13062 3366
rect 13132 3472 13192 3519
rect 13132 3438 13145 3472
rect 13179 3438 13192 3472
rect 13132 3400 13192 3438
rect 13132 3366 13145 3400
rect 13179 3366 13192 3400
rect 13132 3319 13192 3366
rect 13262 3472 13322 3519
rect 13262 3438 13275 3472
rect 13309 3438 13322 3472
rect 13262 3400 13322 3438
rect 13262 3366 13275 3400
rect 13309 3366 13322 3400
rect 13262 3319 13322 3366
rect 13392 3472 13452 3519
rect 13392 3438 13405 3472
rect 13439 3438 13452 3472
rect 13392 3400 13452 3438
rect 13392 3366 13405 3400
rect 13439 3366 13452 3400
rect 13392 3319 13452 3366
rect 13522 3472 13582 3519
rect 13522 3438 13535 3472
rect 13569 3438 13582 3472
rect 13522 3400 13582 3438
rect 13522 3366 13535 3400
rect 13569 3366 13582 3400
rect 13522 3319 13582 3366
rect 13652 3472 13712 3519
rect 13652 3438 13665 3472
rect 13699 3438 13712 3472
rect 13652 3400 13712 3438
rect 13652 3366 13665 3400
rect 13699 3366 13712 3400
rect 13652 3319 13712 3366
rect 13782 3472 13842 3519
rect 13782 3438 13795 3472
rect 13829 3438 13842 3472
rect 13782 3400 13842 3438
rect 13782 3366 13795 3400
rect 13829 3366 13842 3400
rect 13782 3319 13842 3366
rect 13912 3472 13972 3519
rect 13912 3438 13925 3472
rect 13959 3438 13972 3472
rect 13912 3400 13972 3438
rect 13912 3366 13925 3400
rect 13959 3366 13972 3400
rect 13912 3319 13972 3366
rect 14042 3472 14102 3519
rect 14042 3438 14055 3472
rect 14089 3438 14102 3472
rect 14042 3400 14102 3438
rect 14042 3366 14055 3400
rect 14089 3366 14102 3400
rect 14042 3319 14102 3366
rect 14172 3472 14232 3519
rect 14172 3438 14185 3472
rect 14219 3438 14232 3472
rect 14172 3400 14232 3438
rect 14172 3366 14185 3400
rect 14219 3366 14232 3400
rect 14172 3319 14232 3366
rect 14302 3472 14362 3519
rect 14302 3438 14315 3472
rect 14349 3438 14362 3472
rect 14302 3400 14362 3438
rect 14302 3366 14315 3400
rect 14349 3366 14362 3400
rect 14302 3319 14362 3366
rect 14432 3472 14492 3519
rect 14432 3438 14445 3472
rect 14479 3438 14492 3472
rect 14432 3400 14492 3438
rect 14432 3366 14445 3400
rect 14479 3366 14492 3400
rect 14432 3319 14492 3366
rect 14562 3472 14622 3519
rect 14562 3438 14575 3472
rect 14609 3438 14622 3472
rect 14562 3400 14622 3438
rect 14562 3366 14575 3400
rect 14609 3366 14622 3400
rect 14562 3319 14622 3366
rect 14692 3472 14752 3519
rect 14692 3438 14705 3472
rect 14739 3438 14752 3472
rect 14692 3400 14752 3438
rect 14692 3366 14705 3400
rect 14739 3366 14752 3400
rect 14692 3319 14752 3366
rect 14822 3472 14882 3519
rect 14822 3438 14835 3472
rect 14869 3438 14882 3472
rect 14822 3400 14882 3438
rect 14822 3366 14835 3400
rect 14869 3366 14882 3400
rect 14822 3319 14882 3366
rect 14952 3472 15012 3519
rect 14952 3438 14965 3472
rect 14999 3438 15012 3472
rect 14952 3400 15012 3438
rect 14952 3366 14965 3400
rect 14999 3366 15012 3400
rect 14952 3319 15012 3366
rect 15082 3472 15142 3519
rect 15082 3438 15095 3472
rect 15129 3438 15142 3472
rect 15082 3400 15142 3438
rect 15082 3366 15095 3400
rect 15129 3366 15142 3400
rect 15082 3319 15142 3366
rect 24594 3472 24654 3519
rect 24594 3438 24607 3472
rect 24641 3438 24654 3472
rect 24594 3400 24654 3438
rect 24594 3366 24607 3400
rect 24641 3366 24654 3400
rect 24594 3319 24654 3366
rect 24724 3472 24784 3519
rect 24724 3438 24737 3472
rect 24771 3438 24784 3472
rect 24724 3400 24784 3438
rect 24724 3366 24737 3400
rect 24771 3366 24784 3400
rect 24724 3319 24784 3366
rect 24854 3472 24914 3519
rect 24854 3438 24867 3472
rect 24901 3438 24914 3472
rect 24854 3400 24914 3438
rect 24854 3366 24867 3400
rect 24901 3366 24914 3400
rect 24854 3319 24914 3366
rect 24984 3472 25044 3519
rect 24984 3438 24997 3472
rect 25031 3438 25044 3472
rect 24984 3400 25044 3438
rect 24984 3366 24997 3400
rect 25031 3366 25044 3400
rect 24984 3319 25044 3366
rect 25114 3472 25174 3519
rect 25114 3438 25127 3472
rect 25161 3438 25174 3472
rect 25114 3400 25174 3438
rect 25114 3366 25127 3400
rect 25161 3366 25174 3400
rect 25114 3319 25174 3366
rect 25244 3472 25304 3519
rect 25244 3438 25257 3472
rect 25291 3438 25304 3472
rect 25244 3400 25304 3438
rect 25244 3366 25257 3400
rect 25291 3366 25304 3400
rect 25244 3319 25304 3366
rect 25374 3472 25434 3519
rect 25374 3438 25387 3472
rect 25421 3438 25434 3472
rect 25374 3400 25434 3438
rect 25374 3366 25387 3400
rect 25421 3366 25434 3400
rect 25374 3319 25434 3366
rect 25504 3472 25564 3519
rect 25504 3438 25517 3472
rect 25551 3438 25564 3472
rect 25504 3400 25564 3438
rect 25504 3366 25517 3400
rect 25551 3366 25564 3400
rect 25504 3319 25564 3366
rect 25634 3472 25694 3519
rect 25634 3438 25647 3472
rect 25681 3438 25694 3472
rect 25634 3400 25694 3438
rect 25634 3366 25647 3400
rect 25681 3366 25694 3400
rect 25634 3319 25694 3366
rect 25764 3472 25824 3519
rect 25764 3438 25777 3472
rect 25811 3438 25824 3472
rect 25764 3400 25824 3438
rect 25764 3366 25777 3400
rect 25811 3366 25824 3400
rect 25764 3319 25824 3366
rect 25894 3472 25954 3519
rect 25894 3438 25907 3472
rect 25941 3438 25954 3472
rect 25894 3400 25954 3438
rect 25894 3366 25907 3400
rect 25941 3366 25954 3400
rect 25894 3319 25954 3366
rect 26024 3472 26084 3519
rect 26024 3438 26037 3472
rect 26071 3438 26084 3472
rect 26024 3400 26084 3438
rect 26024 3366 26037 3400
rect 26071 3366 26084 3400
rect 26024 3319 26084 3366
rect 26154 3472 26214 3519
rect 26154 3438 26167 3472
rect 26201 3438 26214 3472
rect 26154 3400 26214 3438
rect 26154 3366 26167 3400
rect 26201 3366 26214 3400
rect 26154 3319 26214 3366
rect 26284 3472 26344 3519
rect 26284 3438 26297 3472
rect 26331 3438 26344 3472
rect 26284 3400 26344 3438
rect 26284 3366 26297 3400
rect 26331 3366 26344 3400
rect 26284 3319 26344 3366
rect 26414 3472 26474 3519
rect 26414 3438 26427 3472
rect 26461 3438 26474 3472
rect 26414 3400 26474 3438
rect 26414 3366 26427 3400
rect 26461 3366 26474 3400
rect 26414 3319 26474 3366
rect 26544 3472 26604 3519
rect 26544 3438 26557 3472
rect 26591 3438 26604 3472
rect 26544 3400 26604 3438
rect 26544 3366 26557 3400
rect 26591 3366 26604 3400
rect 26544 3319 26604 3366
rect 26674 3472 26734 3519
rect 26674 3438 26687 3472
rect 26721 3438 26734 3472
rect 26674 3400 26734 3438
rect 26674 3366 26687 3400
rect 26721 3366 26734 3400
rect 26674 3319 26734 3366
rect 13132 2860 13192 2907
rect 13132 2826 13145 2860
rect 13179 2826 13192 2860
rect 13132 2788 13192 2826
rect 13132 2754 13145 2788
rect 13179 2754 13192 2788
rect 13132 2707 13192 2754
rect 13262 2860 13322 2907
rect 13262 2826 13275 2860
rect 13309 2826 13322 2860
rect 13262 2788 13322 2826
rect 13262 2754 13275 2788
rect 13309 2754 13322 2788
rect 13262 2707 13322 2754
rect 13392 2860 13452 2907
rect 13392 2826 13405 2860
rect 13439 2826 13452 2860
rect 13392 2788 13452 2826
rect 13392 2754 13405 2788
rect 13439 2754 13452 2788
rect 13392 2707 13452 2754
rect 13522 2860 13582 2907
rect 13522 2826 13535 2860
rect 13569 2826 13582 2860
rect 13522 2788 13582 2826
rect 13522 2754 13535 2788
rect 13569 2754 13582 2788
rect 13522 2707 13582 2754
rect 13652 2860 13712 2907
rect 13652 2826 13665 2860
rect 13699 2826 13712 2860
rect 13652 2788 13712 2826
rect 13652 2754 13665 2788
rect 13699 2754 13712 2788
rect 13652 2707 13712 2754
rect 13782 2860 13842 2907
rect 13782 2826 13795 2860
rect 13829 2826 13842 2860
rect 13782 2788 13842 2826
rect 13782 2754 13795 2788
rect 13829 2754 13842 2788
rect 13782 2707 13842 2754
rect 13912 2860 13972 2907
rect 13912 2826 13925 2860
rect 13959 2826 13972 2860
rect 13912 2788 13972 2826
rect 13912 2754 13925 2788
rect 13959 2754 13972 2788
rect 13912 2707 13972 2754
rect 14042 2860 14102 2907
rect 14042 2826 14055 2860
rect 14089 2826 14102 2860
rect 14042 2788 14102 2826
rect 14042 2754 14055 2788
rect 14089 2754 14102 2788
rect 14042 2707 14102 2754
rect 14172 2860 14232 2907
rect 14172 2826 14185 2860
rect 14219 2826 14232 2860
rect 14172 2788 14232 2826
rect 14172 2754 14185 2788
rect 14219 2754 14232 2788
rect 14172 2707 14232 2754
rect 14302 2860 14362 2907
rect 14302 2826 14315 2860
rect 14349 2826 14362 2860
rect 14302 2788 14362 2826
rect 14302 2754 14315 2788
rect 14349 2754 14362 2788
rect 14302 2707 14362 2754
rect 14432 2860 14492 2907
rect 14432 2826 14445 2860
rect 14479 2826 14492 2860
rect 14432 2788 14492 2826
rect 14432 2754 14445 2788
rect 14479 2754 14492 2788
rect 14432 2707 14492 2754
rect 14562 2860 14622 2907
rect 14562 2826 14575 2860
rect 14609 2826 14622 2860
rect 14562 2788 14622 2826
rect 14562 2754 14575 2788
rect 14609 2754 14622 2788
rect 14562 2707 14622 2754
rect 14692 2860 14752 2907
rect 14692 2826 14705 2860
rect 14739 2826 14752 2860
rect 14692 2788 14752 2826
rect 14692 2754 14705 2788
rect 14739 2754 14752 2788
rect 14692 2707 14752 2754
rect 14822 2860 14882 2907
rect 14822 2826 14835 2860
rect 14869 2826 14882 2860
rect 14822 2788 14882 2826
rect 14822 2754 14835 2788
rect 14869 2754 14882 2788
rect 14822 2707 14882 2754
rect 14952 2860 15012 2907
rect 14952 2826 14965 2860
rect 14999 2826 15012 2860
rect 14952 2788 15012 2826
rect 14952 2754 14965 2788
rect 14999 2754 15012 2788
rect 14952 2707 15012 2754
rect 15082 2860 15142 2907
rect 15082 2826 15095 2860
rect 15129 2826 15142 2860
rect 15082 2788 15142 2826
rect 15082 2754 15095 2788
rect 15129 2754 15142 2788
rect 15082 2707 15142 2754
rect 15212 2860 15272 2907
rect 15212 2826 15225 2860
rect 15259 2826 15272 2860
rect 15212 2788 15272 2826
rect 15212 2754 15225 2788
rect 15259 2754 15272 2788
rect 15212 2707 15272 2754
rect 15342 2860 15402 2907
rect 15342 2826 15355 2860
rect 15389 2826 15402 2860
rect 15342 2788 15402 2826
rect 15342 2754 15355 2788
rect 15389 2754 15402 2788
rect 15342 2707 15402 2754
rect 15472 2860 15532 2907
rect 15472 2826 15485 2860
rect 15519 2826 15532 2860
rect 15472 2788 15532 2826
rect 15472 2754 15485 2788
rect 15519 2754 15532 2788
rect 15472 2707 15532 2754
rect 24724 2860 24784 2907
rect 24724 2826 24737 2860
rect 24771 2826 24784 2860
rect 24724 2788 24784 2826
rect 24724 2754 24737 2788
rect 24771 2754 24784 2788
rect 24724 2707 24784 2754
rect 24854 2860 24914 2907
rect 24854 2826 24867 2860
rect 24901 2826 24914 2860
rect 24854 2788 24914 2826
rect 24854 2754 24867 2788
rect 24901 2754 24914 2788
rect 24854 2707 24914 2754
rect 24984 2860 25044 2907
rect 24984 2826 24997 2860
rect 25031 2826 25044 2860
rect 24984 2788 25044 2826
rect 24984 2754 24997 2788
rect 25031 2754 25044 2788
rect 24984 2707 25044 2754
rect 25114 2860 25174 2907
rect 25114 2826 25127 2860
rect 25161 2826 25174 2860
rect 25114 2788 25174 2826
rect 25114 2754 25127 2788
rect 25161 2754 25174 2788
rect 25114 2707 25174 2754
rect 25244 2860 25304 2907
rect 25244 2826 25257 2860
rect 25291 2826 25304 2860
rect 25244 2788 25304 2826
rect 25244 2754 25257 2788
rect 25291 2754 25304 2788
rect 25244 2707 25304 2754
rect 25374 2860 25434 2907
rect 25374 2826 25387 2860
rect 25421 2826 25434 2860
rect 25374 2788 25434 2826
rect 25374 2754 25387 2788
rect 25421 2754 25434 2788
rect 25374 2707 25434 2754
rect 25504 2860 25564 2907
rect 25504 2826 25517 2860
rect 25551 2826 25564 2860
rect 25504 2788 25564 2826
rect 25504 2754 25517 2788
rect 25551 2754 25564 2788
rect 25504 2707 25564 2754
rect 25634 2860 25694 2907
rect 25634 2826 25647 2860
rect 25681 2826 25694 2860
rect 25634 2788 25694 2826
rect 25634 2754 25647 2788
rect 25681 2754 25694 2788
rect 25634 2707 25694 2754
rect 25764 2860 25824 2907
rect 25764 2826 25777 2860
rect 25811 2826 25824 2860
rect 25764 2788 25824 2826
rect 25764 2754 25777 2788
rect 25811 2754 25824 2788
rect 25764 2707 25824 2754
rect 25894 2860 25954 2907
rect 25894 2826 25907 2860
rect 25941 2826 25954 2860
rect 25894 2788 25954 2826
rect 25894 2754 25907 2788
rect 25941 2754 25954 2788
rect 25894 2707 25954 2754
rect 26024 2860 26084 2907
rect 26024 2826 26037 2860
rect 26071 2826 26084 2860
rect 26024 2788 26084 2826
rect 26024 2754 26037 2788
rect 26071 2754 26084 2788
rect 26024 2707 26084 2754
rect 26154 2860 26214 2907
rect 26154 2826 26167 2860
rect 26201 2826 26214 2860
rect 26154 2788 26214 2826
rect 26154 2754 26167 2788
rect 26201 2754 26214 2788
rect 26154 2707 26214 2754
rect 26284 2860 26344 2907
rect 26284 2826 26297 2860
rect 26331 2826 26344 2860
rect 26284 2788 26344 2826
rect 26284 2754 26297 2788
rect 26331 2754 26344 2788
rect 26284 2707 26344 2754
rect 26414 2860 26474 2907
rect 26414 2826 26427 2860
rect 26461 2826 26474 2860
rect 26414 2788 26474 2826
rect 26414 2754 26427 2788
rect 26461 2754 26474 2788
rect 26414 2707 26474 2754
rect 26544 2860 26604 2907
rect 26544 2826 26557 2860
rect 26591 2826 26604 2860
rect 26544 2788 26604 2826
rect 26544 2754 26557 2788
rect 26591 2754 26604 2788
rect 26544 2707 26604 2754
rect 26674 2860 26734 2907
rect 26674 2826 26687 2860
rect 26721 2826 26734 2860
rect 26674 2788 26734 2826
rect 26674 2754 26687 2788
rect 26721 2754 26734 2788
rect 26674 2707 26734 2754
rect 26804 2860 26864 2907
rect 26804 2826 26817 2860
rect 26851 2826 26864 2860
rect 26804 2788 26864 2826
rect 26804 2754 26817 2788
rect 26851 2754 26864 2788
rect 26804 2707 26864 2754
rect 26934 2860 26994 2907
rect 26934 2826 26947 2860
rect 26981 2826 26994 2860
rect 26934 2788 26994 2826
rect 26934 2754 26947 2788
rect 26981 2754 26994 2788
rect 26934 2707 26994 2754
rect 27064 2860 27124 2907
rect 27064 2826 27077 2860
rect 27111 2826 27124 2860
rect 27064 2788 27124 2826
rect 27064 2754 27077 2788
rect 27111 2754 27124 2788
rect 27064 2707 27124 2754
rect 13132 2512 13192 2559
rect 13132 2478 13145 2512
rect 13179 2478 13192 2512
rect 13132 2440 13192 2478
rect 13132 2406 13145 2440
rect 13179 2406 13192 2440
rect 13132 2359 13192 2406
rect 13262 2512 13322 2559
rect 13262 2478 13275 2512
rect 13309 2478 13322 2512
rect 13262 2440 13322 2478
rect 13262 2406 13275 2440
rect 13309 2406 13322 2440
rect 13262 2359 13322 2406
rect 13392 2512 13452 2559
rect 13392 2478 13405 2512
rect 13439 2478 13452 2512
rect 13392 2440 13452 2478
rect 13392 2406 13405 2440
rect 13439 2406 13452 2440
rect 13392 2359 13452 2406
rect 13522 2512 13582 2559
rect 13522 2478 13535 2512
rect 13569 2478 13582 2512
rect 13522 2440 13582 2478
rect 13522 2406 13535 2440
rect 13569 2406 13582 2440
rect 13522 2359 13582 2406
rect 13652 2512 13712 2559
rect 13652 2478 13665 2512
rect 13699 2478 13712 2512
rect 13652 2440 13712 2478
rect 13652 2406 13665 2440
rect 13699 2406 13712 2440
rect 13652 2359 13712 2406
rect 13782 2512 13842 2559
rect 13782 2478 13795 2512
rect 13829 2478 13842 2512
rect 13782 2440 13842 2478
rect 13782 2406 13795 2440
rect 13829 2406 13842 2440
rect 13782 2359 13842 2406
rect 13912 2512 13972 2559
rect 13912 2478 13925 2512
rect 13959 2478 13972 2512
rect 13912 2440 13972 2478
rect 13912 2406 13925 2440
rect 13959 2406 13972 2440
rect 13912 2359 13972 2406
rect 14042 2512 14102 2559
rect 14042 2478 14055 2512
rect 14089 2478 14102 2512
rect 14042 2440 14102 2478
rect 14042 2406 14055 2440
rect 14089 2406 14102 2440
rect 14042 2359 14102 2406
rect 14172 2512 14232 2559
rect 14172 2478 14185 2512
rect 14219 2478 14232 2512
rect 14172 2440 14232 2478
rect 14172 2406 14185 2440
rect 14219 2406 14232 2440
rect 14172 2359 14232 2406
rect 14302 2512 14362 2559
rect 14302 2478 14315 2512
rect 14349 2478 14362 2512
rect 14302 2440 14362 2478
rect 14302 2406 14315 2440
rect 14349 2406 14362 2440
rect 14302 2359 14362 2406
rect 14432 2512 14492 2559
rect 14432 2478 14445 2512
rect 14479 2478 14492 2512
rect 14432 2440 14492 2478
rect 14432 2406 14445 2440
rect 14479 2406 14492 2440
rect 14432 2359 14492 2406
rect 14562 2512 14622 2559
rect 14562 2478 14575 2512
rect 14609 2478 14622 2512
rect 14562 2440 14622 2478
rect 14562 2406 14575 2440
rect 14609 2406 14622 2440
rect 14562 2359 14622 2406
rect 14692 2512 14752 2559
rect 14692 2478 14705 2512
rect 14739 2478 14752 2512
rect 14692 2440 14752 2478
rect 14692 2406 14705 2440
rect 14739 2406 14752 2440
rect 14692 2359 14752 2406
rect 14822 2512 14882 2559
rect 14822 2478 14835 2512
rect 14869 2478 14882 2512
rect 14822 2440 14882 2478
rect 14822 2406 14835 2440
rect 14869 2406 14882 2440
rect 14822 2359 14882 2406
rect 14952 2512 15012 2559
rect 14952 2478 14965 2512
rect 14999 2478 15012 2512
rect 14952 2440 15012 2478
rect 14952 2406 14965 2440
rect 14999 2406 15012 2440
rect 14952 2359 15012 2406
rect 15082 2512 15142 2559
rect 15082 2478 15095 2512
rect 15129 2478 15142 2512
rect 15082 2440 15142 2478
rect 15082 2406 15095 2440
rect 15129 2406 15142 2440
rect 15082 2359 15142 2406
rect 15212 2512 15272 2559
rect 15212 2478 15225 2512
rect 15259 2478 15272 2512
rect 15212 2440 15272 2478
rect 15212 2406 15225 2440
rect 15259 2406 15272 2440
rect 15212 2359 15272 2406
rect 15342 2512 15402 2559
rect 15342 2478 15355 2512
rect 15389 2478 15402 2512
rect 15342 2440 15402 2478
rect 15342 2406 15355 2440
rect 15389 2406 15402 2440
rect 15342 2359 15402 2406
rect 24724 2512 24784 2559
rect 24724 2478 24737 2512
rect 24771 2478 24784 2512
rect 24724 2440 24784 2478
rect 24724 2406 24737 2440
rect 24771 2406 24784 2440
rect 24724 2359 24784 2406
rect 24854 2512 24914 2559
rect 24854 2478 24867 2512
rect 24901 2478 24914 2512
rect 24854 2440 24914 2478
rect 24854 2406 24867 2440
rect 24901 2406 24914 2440
rect 24854 2359 24914 2406
rect 24984 2512 25044 2559
rect 24984 2478 24997 2512
rect 25031 2478 25044 2512
rect 24984 2440 25044 2478
rect 24984 2406 24997 2440
rect 25031 2406 25044 2440
rect 24984 2359 25044 2406
rect 25114 2512 25174 2559
rect 25114 2478 25127 2512
rect 25161 2478 25174 2512
rect 25114 2440 25174 2478
rect 25114 2406 25127 2440
rect 25161 2406 25174 2440
rect 25114 2359 25174 2406
rect 25244 2512 25304 2559
rect 25244 2478 25257 2512
rect 25291 2478 25304 2512
rect 25244 2440 25304 2478
rect 25244 2406 25257 2440
rect 25291 2406 25304 2440
rect 25244 2359 25304 2406
rect 25374 2512 25434 2559
rect 25374 2478 25387 2512
rect 25421 2478 25434 2512
rect 25374 2440 25434 2478
rect 25374 2406 25387 2440
rect 25421 2406 25434 2440
rect 25374 2359 25434 2406
rect 25504 2512 25564 2559
rect 25504 2478 25517 2512
rect 25551 2478 25564 2512
rect 25504 2440 25564 2478
rect 25504 2406 25517 2440
rect 25551 2406 25564 2440
rect 25504 2359 25564 2406
rect 25634 2512 25694 2559
rect 25634 2478 25647 2512
rect 25681 2478 25694 2512
rect 25634 2440 25694 2478
rect 25634 2406 25647 2440
rect 25681 2406 25694 2440
rect 25634 2359 25694 2406
rect 25764 2512 25824 2559
rect 25764 2478 25777 2512
rect 25811 2478 25824 2512
rect 25764 2440 25824 2478
rect 25764 2406 25777 2440
rect 25811 2406 25824 2440
rect 25764 2359 25824 2406
rect 25894 2512 25954 2559
rect 25894 2478 25907 2512
rect 25941 2478 25954 2512
rect 25894 2440 25954 2478
rect 25894 2406 25907 2440
rect 25941 2406 25954 2440
rect 25894 2359 25954 2406
rect 26024 2512 26084 2559
rect 26024 2478 26037 2512
rect 26071 2478 26084 2512
rect 26024 2440 26084 2478
rect 26024 2406 26037 2440
rect 26071 2406 26084 2440
rect 26024 2359 26084 2406
rect 26154 2512 26214 2559
rect 26154 2478 26167 2512
rect 26201 2478 26214 2512
rect 26154 2440 26214 2478
rect 26154 2406 26167 2440
rect 26201 2406 26214 2440
rect 26154 2359 26214 2406
rect 26284 2512 26344 2559
rect 26284 2478 26297 2512
rect 26331 2478 26344 2512
rect 26284 2440 26344 2478
rect 26284 2406 26297 2440
rect 26331 2406 26344 2440
rect 26284 2359 26344 2406
rect 26414 2512 26474 2559
rect 26414 2478 26427 2512
rect 26461 2478 26474 2512
rect 26414 2440 26474 2478
rect 26414 2406 26427 2440
rect 26461 2406 26474 2440
rect 26414 2359 26474 2406
rect 26544 2512 26604 2559
rect 26544 2478 26557 2512
rect 26591 2478 26604 2512
rect 26544 2440 26604 2478
rect 26544 2406 26557 2440
rect 26591 2406 26604 2440
rect 26544 2359 26604 2406
rect 26674 2512 26734 2559
rect 26674 2478 26687 2512
rect 26721 2478 26734 2512
rect 26674 2440 26734 2478
rect 26674 2406 26687 2440
rect 26721 2406 26734 2440
rect 26674 2359 26734 2406
rect 26804 2512 26864 2559
rect 26804 2478 26817 2512
rect 26851 2478 26864 2512
rect 26804 2440 26864 2478
rect 26804 2406 26817 2440
rect 26851 2406 26864 2440
rect 26804 2359 26864 2406
rect 26934 2512 26994 2559
rect 26934 2478 26947 2512
rect 26981 2478 26994 2512
rect 26934 2440 26994 2478
rect 26934 2406 26947 2440
rect 26981 2406 26994 2440
rect 26934 2359 26994 2406
<< pdiff >>
rect 13002 5224 13062 5263
rect 13002 5190 13015 5224
rect 13049 5190 13062 5224
rect 13002 5152 13062 5190
rect 13002 5118 13015 5152
rect 13049 5118 13062 5152
rect 13002 5080 13062 5118
rect 13002 5046 13015 5080
rect 13049 5046 13062 5080
rect 13002 5008 13062 5046
rect 13002 4974 13015 5008
rect 13049 4974 13062 5008
rect 13002 4936 13062 4974
rect 13002 4902 13015 4936
rect 13049 4902 13062 4936
rect 13002 4863 13062 4902
rect 13132 5224 13192 5263
rect 13132 5190 13145 5224
rect 13179 5190 13192 5224
rect 13132 5152 13192 5190
rect 13132 5118 13145 5152
rect 13179 5118 13192 5152
rect 13132 5080 13192 5118
rect 13132 5046 13145 5080
rect 13179 5046 13192 5080
rect 13132 5008 13192 5046
rect 13132 4974 13145 5008
rect 13179 4974 13192 5008
rect 13132 4936 13192 4974
rect 13132 4902 13145 4936
rect 13179 4902 13192 4936
rect 13132 4863 13192 4902
rect 13262 5224 13322 5263
rect 13262 5190 13275 5224
rect 13309 5190 13322 5224
rect 13262 5152 13322 5190
rect 13262 5118 13275 5152
rect 13309 5118 13322 5152
rect 13262 5080 13322 5118
rect 13262 5046 13275 5080
rect 13309 5046 13322 5080
rect 13262 5008 13322 5046
rect 13262 4974 13275 5008
rect 13309 4974 13322 5008
rect 13262 4936 13322 4974
rect 13262 4902 13275 4936
rect 13309 4902 13322 4936
rect 13262 4863 13322 4902
rect 13392 5224 13452 5263
rect 13392 5190 13405 5224
rect 13439 5190 13452 5224
rect 13392 5152 13452 5190
rect 13392 5118 13405 5152
rect 13439 5118 13452 5152
rect 13392 5080 13452 5118
rect 13392 5046 13405 5080
rect 13439 5046 13452 5080
rect 13392 5008 13452 5046
rect 13392 4974 13405 5008
rect 13439 4974 13452 5008
rect 13392 4936 13452 4974
rect 13392 4902 13405 4936
rect 13439 4902 13452 4936
rect 13392 4863 13452 4902
rect 13522 5224 13582 5263
rect 13522 5190 13535 5224
rect 13569 5190 13582 5224
rect 13522 5152 13582 5190
rect 13522 5118 13535 5152
rect 13569 5118 13582 5152
rect 13522 5080 13582 5118
rect 13522 5046 13535 5080
rect 13569 5046 13582 5080
rect 13522 5008 13582 5046
rect 13522 4974 13535 5008
rect 13569 4974 13582 5008
rect 13522 4936 13582 4974
rect 13522 4902 13535 4936
rect 13569 4902 13582 4936
rect 13522 4863 13582 4902
rect 13652 5224 13712 5263
rect 13652 5190 13665 5224
rect 13699 5190 13712 5224
rect 13652 5152 13712 5190
rect 13652 5118 13665 5152
rect 13699 5118 13712 5152
rect 13652 5080 13712 5118
rect 13652 5046 13665 5080
rect 13699 5046 13712 5080
rect 13652 5008 13712 5046
rect 13652 4974 13665 5008
rect 13699 4974 13712 5008
rect 13652 4936 13712 4974
rect 13652 4902 13665 4936
rect 13699 4902 13712 4936
rect 13652 4863 13712 4902
rect 13782 5224 13842 5263
rect 13782 5190 13795 5224
rect 13829 5190 13842 5224
rect 13782 5152 13842 5190
rect 13782 5118 13795 5152
rect 13829 5118 13842 5152
rect 13782 5080 13842 5118
rect 13782 5046 13795 5080
rect 13829 5046 13842 5080
rect 13782 5008 13842 5046
rect 13782 4974 13795 5008
rect 13829 4974 13842 5008
rect 13782 4936 13842 4974
rect 13782 4902 13795 4936
rect 13829 4902 13842 4936
rect 13782 4863 13842 4902
rect 13912 5224 13972 5263
rect 13912 5190 13925 5224
rect 13959 5190 13972 5224
rect 13912 5152 13972 5190
rect 13912 5118 13925 5152
rect 13959 5118 13972 5152
rect 13912 5080 13972 5118
rect 13912 5046 13925 5080
rect 13959 5046 13972 5080
rect 13912 5008 13972 5046
rect 13912 4974 13925 5008
rect 13959 4974 13972 5008
rect 13912 4936 13972 4974
rect 13912 4902 13925 4936
rect 13959 4902 13972 4936
rect 13912 4863 13972 4902
rect 14042 5224 14102 5263
rect 14042 5190 14055 5224
rect 14089 5190 14102 5224
rect 14042 5152 14102 5190
rect 14042 5118 14055 5152
rect 14089 5118 14102 5152
rect 14042 5080 14102 5118
rect 14042 5046 14055 5080
rect 14089 5046 14102 5080
rect 14042 5008 14102 5046
rect 14042 4974 14055 5008
rect 14089 4974 14102 5008
rect 14042 4936 14102 4974
rect 14042 4902 14055 4936
rect 14089 4902 14102 4936
rect 14042 4863 14102 4902
rect 14172 5224 14232 5263
rect 14172 5190 14185 5224
rect 14219 5190 14232 5224
rect 14172 5152 14232 5190
rect 14172 5118 14185 5152
rect 14219 5118 14232 5152
rect 14172 5080 14232 5118
rect 14172 5046 14185 5080
rect 14219 5046 14232 5080
rect 14172 5008 14232 5046
rect 14172 4974 14185 5008
rect 14219 4974 14232 5008
rect 14172 4936 14232 4974
rect 14172 4902 14185 4936
rect 14219 4902 14232 4936
rect 14172 4863 14232 4902
rect 14302 5224 14362 5263
rect 14302 5190 14315 5224
rect 14349 5190 14362 5224
rect 14302 5152 14362 5190
rect 14302 5118 14315 5152
rect 14349 5118 14362 5152
rect 14302 5080 14362 5118
rect 14302 5046 14315 5080
rect 14349 5046 14362 5080
rect 14302 5008 14362 5046
rect 14302 4974 14315 5008
rect 14349 4974 14362 5008
rect 14302 4936 14362 4974
rect 14302 4902 14315 4936
rect 14349 4902 14362 4936
rect 14302 4863 14362 4902
rect 14432 5224 14492 5263
rect 14432 5190 14445 5224
rect 14479 5190 14492 5224
rect 14432 5152 14492 5190
rect 14432 5118 14445 5152
rect 14479 5118 14492 5152
rect 14432 5080 14492 5118
rect 14432 5046 14445 5080
rect 14479 5046 14492 5080
rect 14432 5008 14492 5046
rect 14432 4974 14445 5008
rect 14479 4974 14492 5008
rect 14432 4936 14492 4974
rect 14432 4902 14445 4936
rect 14479 4902 14492 4936
rect 14432 4863 14492 4902
rect 14562 5224 14622 5263
rect 14562 5190 14575 5224
rect 14609 5190 14622 5224
rect 14562 5152 14622 5190
rect 14562 5118 14575 5152
rect 14609 5118 14622 5152
rect 14562 5080 14622 5118
rect 14562 5046 14575 5080
rect 14609 5046 14622 5080
rect 14562 5008 14622 5046
rect 14562 4974 14575 5008
rect 14609 4974 14622 5008
rect 14562 4936 14622 4974
rect 14562 4902 14575 4936
rect 14609 4902 14622 4936
rect 14562 4863 14622 4902
rect 14692 5224 14752 5263
rect 14692 5190 14705 5224
rect 14739 5190 14752 5224
rect 14692 5152 14752 5190
rect 14692 5118 14705 5152
rect 14739 5118 14752 5152
rect 14692 5080 14752 5118
rect 14692 5046 14705 5080
rect 14739 5046 14752 5080
rect 14692 5008 14752 5046
rect 14692 4974 14705 5008
rect 14739 4974 14752 5008
rect 14692 4936 14752 4974
rect 14692 4902 14705 4936
rect 14739 4902 14752 4936
rect 14692 4863 14752 4902
rect 14822 5224 14882 5263
rect 14822 5190 14835 5224
rect 14869 5190 14882 5224
rect 14822 5152 14882 5190
rect 14822 5118 14835 5152
rect 14869 5118 14882 5152
rect 14822 5080 14882 5118
rect 14822 5046 14835 5080
rect 14869 5046 14882 5080
rect 14822 5008 14882 5046
rect 14822 4974 14835 5008
rect 14869 4974 14882 5008
rect 14822 4936 14882 4974
rect 14822 4902 14835 4936
rect 14869 4902 14882 4936
rect 14822 4863 14882 4902
rect 14952 5224 15012 5263
rect 14952 5190 14965 5224
rect 14999 5190 15012 5224
rect 14952 5152 15012 5190
rect 14952 5118 14965 5152
rect 14999 5118 15012 5152
rect 14952 5080 15012 5118
rect 14952 5046 14965 5080
rect 14999 5046 15012 5080
rect 14952 5008 15012 5046
rect 14952 4974 14965 5008
rect 14999 4974 15012 5008
rect 14952 4936 15012 4974
rect 14952 4902 14965 4936
rect 14999 4902 15012 4936
rect 14952 4863 15012 4902
rect 15082 5224 15142 5263
rect 15082 5190 15095 5224
rect 15129 5190 15142 5224
rect 15082 5152 15142 5190
rect 15082 5118 15095 5152
rect 15129 5118 15142 5152
rect 15082 5080 15142 5118
rect 15082 5046 15095 5080
rect 15129 5046 15142 5080
rect 15082 5008 15142 5046
rect 15082 4974 15095 5008
rect 15129 4974 15142 5008
rect 15082 4936 15142 4974
rect 15082 4902 15095 4936
rect 15129 4902 15142 4936
rect 24594 5224 24654 5263
rect 24594 5190 24607 5224
rect 24641 5190 24654 5224
rect 24594 5152 24654 5190
rect 24594 5118 24607 5152
rect 24641 5118 24654 5152
rect 24594 5080 24654 5118
rect 24594 5046 24607 5080
rect 24641 5046 24654 5080
rect 24594 5008 24654 5046
rect 24594 4974 24607 5008
rect 24641 4974 24654 5008
rect 24594 4936 24654 4974
rect 15082 4863 15142 4902
rect 24594 4902 24607 4936
rect 24641 4902 24654 4936
rect 24594 4863 24654 4902
rect 24724 5224 24784 5263
rect 24724 5190 24737 5224
rect 24771 5190 24784 5224
rect 24724 5152 24784 5190
rect 24724 5118 24737 5152
rect 24771 5118 24784 5152
rect 24724 5080 24784 5118
rect 24724 5046 24737 5080
rect 24771 5046 24784 5080
rect 24724 5008 24784 5046
rect 24724 4974 24737 5008
rect 24771 4974 24784 5008
rect 24724 4936 24784 4974
rect 24724 4902 24737 4936
rect 24771 4902 24784 4936
rect 24724 4863 24784 4902
rect 24854 5224 24914 5263
rect 24854 5190 24867 5224
rect 24901 5190 24914 5224
rect 24854 5152 24914 5190
rect 24854 5118 24867 5152
rect 24901 5118 24914 5152
rect 24854 5080 24914 5118
rect 24854 5046 24867 5080
rect 24901 5046 24914 5080
rect 24854 5008 24914 5046
rect 24854 4974 24867 5008
rect 24901 4974 24914 5008
rect 24854 4936 24914 4974
rect 24854 4902 24867 4936
rect 24901 4902 24914 4936
rect 24854 4863 24914 4902
rect 24984 5224 25044 5263
rect 24984 5190 24997 5224
rect 25031 5190 25044 5224
rect 24984 5152 25044 5190
rect 24984 5118 24997 5152
rect 25031 5118 25044 5152
rect 24984 5080 25044 5118
rect 24984 5046 24997 5080
rect 25031 5046 25044 5080
rect 24984 5008 25044 5046
rect 24984 4974 24997 5008
rect 25031 4974 25044 5008
rect 24984 4936 25044 4974
rect 24984 4902 24997 4936
rect 25031 4902 25044 4936
rect 24984 4863 25044 4902
rect 25114 5224 25174 5263
rect 25114 5190 25127 5224
rect 25161 5190 25174 5224
rect 25114 5152 25174 5190
rect 25114 5118 25127 5152
rect 25161 5118 25174 5152
rect 25114 5080 25174 5118
rect 25114 5046 25127 5080
rect 25161 5046 25174 5080
rect 25114 5008 25174 5046
rect 25114 4974 25127 5008
rect 25161 4974 25174 5008
rect 25114 4936 25174 4974
rect 25114 4902 25127 4936
rect 25161 4902 25174 4936
rect 25114 4863 25174 4902
rect 25244 5224 25304 5263
rect 25244 5190 25257 5224
rect 25291 5190 25304 5224
rect 25244 5152 25304 5190
rect 25244 5118 25257 5152
rect 25291 5118 25304 5152
rect 25244 5080 25304 5118
rect 25244 5046 25257 5080
rect 25291 5046 25304 5080
rect 25244 5008 25304 5046
rect 25244 4974 25257 5008
rect 25291 4974 25304 5008
rect 25244 4936 25304 4974
rect 25244 4902 25257 4936
rect 25291 4902 25304 4936
rect 25244 4863 25304 4902
rect 25374 5224 25434 5263
rect 25374 5190 25387 5224
rect 25421 5190 25434 5224
rect 25374 5152 25434 5190
rect 25374 5118 25387 5152
rect 25421 5118 25434 5152
rect 25374 5080 25434 5118
rect 25374 5046 25387 5080
rect 25421 5046 25434 5080
rect 25374 5008 25434 5046
rect 25374 4974 25387 5008
rect 25421 4974 25434 5008
rect 25374 4936 25434 4974
rect 25374 4902 25387 4936
rect 25421 4902 25434 4936
rect 25374 4863 25434 4902
rect 25504 5224 25564 5263
rect 25504 5190 25517 5224
rect 25551 5190 25564 5224
rect 25504 5152 25564 5190
rect 25504 5118 25517 5152
rect 25551 5118 25564 5152
rect 25504 5080 25564 5118
rect 25504 5046 25517 5080
rect 25551 5046 25564 5080
rect 25504 5008 25564 5046
rect 25504 4974 25517 5008
rect 25551 4974 25564 5008
rect 25504 4936 25564 4974
rect 25504 4902 25517 4936
rect 25551 4902 25564 4936
rect 25504 4863 25564 4902
rect 25634 5224 25694 5263
rect 25634 5190 25647 5224
rect 25681 5190 25694 5224
rect 25634 5152 25694 5190
rect 25634 5118 25647 5152
rect 25681 5118 25694 5152
rect 25634 5080 25694 5118
rect 25634 5046 25647 5080
rect 25681 5046 25694 5080
rect 25634 5008 25694 5046
rect 25634 4974 25647 5008
rect 25681 4974 25694 5008
rect 25634 4936 25694 4974
rect 25634 4902 25647 4936
rect 25681 4902 25694 4936
rect 25634 4863 25694 4902
rect 25764 5224 25824 5263
rect 25764 5190 25777 5224
rect 25811 5190 25824 5224
rect 25764 5152 25824 5190
rect 25764 5118 25777 5152
rect 25811 5118 25824 5152
rect 25764 5080 25824 5118
rect 25764 5046 25777 5080
rect 25811 5046 25824 5080
rect 25764 5008 25824 5046
rect 25764 4974 25777 5008
rect 25811 4974 25824 5008
rect 25764 4936 25824 4974
rect 25764 4902 25777 4936
rect 25811 4902 25824 4936
rect 25764 4863 25824 4902
rect 25894 5224 25954 5263
rect 25894 5190 25907 5224
rect 25941 5190 25954 5224
rect 25894 5152 25954 5190
rect 25894 5118 25907 5152
rect 25941 5118 25954 5152
rect 25894 5080 25954 5118
rect 25894 5046 25907 5080
rect 25941 5046 25954 5080
rect 25894 5008 25954 5046
rect 25894 4974 25907 5008
rect 25941 4974 25954 5008
rect 25894 4936 25954 4974
rect 25894 4902 25907 4936
rect 25941 4902 25954 4936
rect 25894 4863 25954 4902
rect 26024 5224 26084 5263
rect 26024 5190 26037 5224
rect 26071 5190 26084 5224
rect 26024 5152 26084 5190
rect 26024 5118 26037 5152
rect 26071 5118 26084 5152
rect 26024 5080 26084 5118
rect 26024 5046 26037 5080
rect 26071 5046 26084 5080
rect 26024 5008 26084 5046
rect 26024 4974 26037 5008
rect 26071 4974 26084 5008
rect 26024 4936 26084 4974
rect 26024 4902 26037 4936
rect 26071 4902 26084 4936
rect 26024 4863 26084 4902
rect 26154 5224 26214 5263
rect 26154 5190 26167 5224
rect 26201 5190 26214 5224
rect 26154 5152 26214 5190
rect 26154 5118 26167 5152
rect 26201 5118 26214 5152
rect 26154 5080 26214 5118
rect 26154 5046 26167 5080
rect 26201 5046 26214 5080
rect 26154 5008 26214 5046
rect 26154 4974 26167 5008
rect 26201 4974 26214 5008
rect 26154 4936 26214 4974
rect 26154 4902 26167 4936
rect 26201 4902 26214 4936
rect 26154 4863 26214 4902
rect 26284 5224 26344 5263
rect 26284 5190 26297 5224
rect 26331 5190 26344 5224
rect 26284 5152 26344 5190
rect 26284 5118 26297 5152
rect 26331 5118 26344 5152
rect 26284 5080 26344 5118
rect 26284 5046 26297 5080
rect 26331 5046 26344 5080
rect 26284 5008 26344 5046
rect 26284 4974 26297 5008
rect 26331 4974 26344 5008
rect 26284 4936 26344 4974
rect 26284 4902 26297 4936
rect 26331 4902 26344 4936
rect 26284 4863 26344 4902
rect 26414 5224 26474 5263
rect 26414 5190 26427 5224
rect 26461 5190 26474 5224
rect 26414 5152 26474 5190
rect 26414 5118 26427 5152
rect 26461 5118 26474 5152
rect 26414 5080 26474 5118
rect 26414 5046 26427 5080
rect 26461 5046 26474 5080
rect 26414 5008 26474 5046
rect 26414 4974 26427 5008
rect 26461 4974 26474 5008
rect 26414 4936 26474 4974
rect 26414 4902 26427 4936
rect 26461 4902 26474 4936
rect 26414 4863 26474 4902
rect 26544 5224 26604 5263
rect 26544 5190 26557 5224
rect 26591 5190 26604 5224
rect 26544 5152 26604 5190
rect 26544 5118 26557 5152
rect 26591 5118 26604 5152
rect 26544 5080 26604 5118
rect 26544 5046 26557 5080
rect 26591 5046 26604 5080
rect 26544 5008 26604 5046
rect 26544 4974 26557 5008
rect 26591 4974 26604 5008
rect 26544 4936 26604 4974
rect 26544 4902 26557 4936
rect 26591 4902 26604 4936
rect 26544 4863 26604 4902
rect 26674 5224 26734 5263
rect 26674 5190 26687 5224
rect 26721 5190 26734 5224
rect 26674 5152 26734 5190
rect 26674 5118 26687 5152
rect 26721 5118 26734 5152
rect 26674 5080 26734 5118
rect 26674 5046 26687 5080
rect 26721 5046 26734 5080
rect 26674 5008 26734 5046
rect 26674 4974 26687 5008
rect 26721 4974 26734 5008
rect 26674 4936 26734 4974
rect 26674 4902 26687 4936
rect 26721 4902 26734 4936
rect 26674 4863 26734 4902
rect 13262 4676 13322 4715
rect 13262 4642 13275 4676
rect 13309 4642 13322 4676
rect 13262 4604 13322 4642
rect 13262 4570 13275 4604
rect 13309 4570 13322 4604
rect 13262 4532 13322 4570
rect 13262 4498 13275 4532
rect 13309 4498 13322 4532
rect 13262 4460 13322 4498
rect 13262 4426 13275 4460
rect 13309 4426 13322 4460
rect 13262 4388 13322 4426
rect 13262 4354 13275 4388
rect 13309 4354 13322 4388
rect 13262 4315 13322 4354
rect 13392 4676 13452 4715
rect 13392 4642 13405 4676
rect 13439 4642 13452 4676
rect 13392 4604 13452 4642
rect 13392 4570 13405 4604
rect 13439 4570 13452 4604
rect 13392 4532 13452 4570
rect 13392 4498 13405 4532
rect 13439 4498 13452 4532
rect 13392 4460 13452 4498
rect 13392 4426 13405 4460
rect 13439 4426 13452 4460
rect 13392 4388 13452 4426
rect 13392 4354 13405 4388
rect 13439 4354 13452 4388
rect 13392 4315 13452 4354
rect 13652 4676 13712 4715
rect 13652 4642 13665 4676
rect 13699 4642 13712 4676
rect 13652 4604 13712 4642
rect 13652 4570 13665 4604
rect 13699 4570 13712 4604
rect 13652 4532 13712 4570
rect 13652 4498 13665 4532
rect 13699 4498 13712 4532
rect 13652 4460 13712 4498
rect 13652 4426 13665 4460
rect 13699 4426 13712 4460
rect 13652 4388 13712 4426
rect 13652 4354 13665 4388
rect 13699 4354 13712 4388
rect 13652 4315 13712 4354
rect 13782 4676 13842 4715
rect 13782 4642 13795 4676
rect 13829 4642 13842 4676
rect 13782 4604 13842 4642
rect 13782 4570 13795 4604
rect 13829 4570 13842 4604
rect 13782 4532 13842 4570
rect 13782 4498 13795 4532
rect 13829 4498 13842 4532
rect 13782 4460 13842 4498
rect 13782 4426 13795 4460
rect 13829 4426 13842 4460
rect 13782 4388 13842 4426
rect 13782 4354 13795 4388
rect 13829 4354 13842 4388
rect 13782 4315 13842 4354
rect 14042 4676 14102 4715
rect 14042 4642 14055 4676
rect 14089 4642 14102 4676
rect 14042 4604 14102 4642
rect 14042 4570 14055 4604
rect 14089 4570 14102 4604
rect 14042 4532 14102 4570
rect 14042 4498 14055 4532
rect 14089 4498 14102 4532
rect 14042 4460 14102 4498
rect 14042 4426 14055 4460
rect 14089 4426 14102 4460
rect 14042 4388 14102 4426
rect 14042 4354 14055 4388
rect 14089 4354 14102 4388
rect 14042 4315 14102 4354
rect 14172 4676 14232 4715
rect 14172 4642 14185 4676
rect 14219 4642 14232 4676
rect 14172 4604 14232 4642
rect 14172 4570 14185 4604
rect 14219 4570 14232 4604
rect 14172 4532 14232 4570
rect 14172 4498 14185 4532
rect 14219 4498 14232 4532
rect 14172 4460 14232 4498
rect 14172 4426 14185 4460
rect 14219 4426 14232 4460
rect 14172 4388 14232 4426
rect 14172 4354 14185 4388
rect 14219 4354 14232 4388
rect 14172 4315 14232 4354
rect 14432 4676 14492 4715
rect 14432 4642 14445 4676
rect 14479 4642 14492 4676
rect 14432 4604 14492 4642
rect 14432 4570 14445 4604
rect 14479 4570 14492 4604
rect 14432 4532 14492 4570
rect 14432 4498 14445 4532
rect 14479 4498 14492 4532
rect 14432 4460 14492 4498
rect 14432 4426 14445 4460
rect 14479 4426 14492 4460
rect 14432 4388 14492 4426
rect 14432 4354 14445 4388
rect 14479 4354 14492 4388
rect 14432 4315 14492 4354
rect 14562 4676 14622 4715
rect 14562 4642 14575 4676
rect 14609 4642 14622 4676
rect 14562 4604 14622 4642
rect 14562 4570 14575 4604
rect 14609 4570 14622 4604
rect 14562 4532 14622 4570
rect 14562 4498 14575 4532
rect 14609 4498 14622 4532
rect 14562 4460 14622 4498
rect 14562 4426 14575 4460
rect 14609 4426 14622 4460
rect 14562 4388 14622 4426
rect 14562 4354 14575 4388
rect 14609 4354 14622 4388
rect 14562 4315 14622 4354
rect 14822 4676 14882 4715
rect 14822 4642 14835 4676
rect 14869 4642 14882 4676
rect 14822 4604 14882 4642
rect 14822 4570 14835 4604
rect 14869 4570 14882 4604
rect 14822 4532 14882 4570
rect 14822 4498 14835 4532
rect 14869 4498 14882 4532
rect 14822 4460 14882 4498
rect 14822 4426 14835 4460
rect 14869 4426 14882 4460
rect 14822 4388 14882 4426
rect 14822 4354 14835 4388
rect 14869 4354 14882 4388
rect 14822 4315 14882 4354
rect 14952 4676 15012 4715
rect 14952 4642 14965 4676
rect 14999 4642 15012 4676
rect 14952 4604 15012 4642
rect 14952 4570 14965 4604
rect 14999 4570 15012 4604
rect 14952 4532 15012 4570
rect 14952 4498 14965 4532
rect 14999 4498 15012 4532
rect 14952 4460 15012 4498
rect 14952 4426 14965 4460
rect 14999 4426 15012 4460
rect 14952 4388 15012 4426
rect 14952 4354 14965 4388
rect 14999 4354 15012 4388
rect 14952 4315 15012 4354
rect 15196 4676 15256 4715
rect 15196 4642 15209 4676
rect 15243 4642 15256 4676
rect 15196 4604 15256 4642
rect 15196 4570 15209 4604
rect 15243 4570 15256 4604
rect 15196 4532 15256 4570
rect 15196 4498 15209 4532
rect 15243 4498 15256 4532
rect 15196 4460 15256 4498
rect 15196 4426 15209 4460
rect 15243 4426 15256 4460
rect 15196 4388 15256 4426
rect 15196 4354 15209 4388
rect 15243 4354 15256 4388
rect 15196 4315 15256 4354
rect 15286 4676 15346 4715
rect 15286 4642 15299 4676
rect 15333 4642 15346 4676
rect 15286 4604 15346 4642
rect 15286 4570 15299 4604
rect 15333 4570 15346 4604
rect 15286 4532 15346 4570
rect 15286 4498 15299 4532
rect 15333 4498 15346 4532
rect 15286 4460 15346 4498
rect 15286 4426 15299 4460
rect 15333 4426 15346 4460
rect 15286 4388 15346 4426
rect 15286 4354 15299 4388
rect 15333 4354 15346 4388
rect 15286 4315 15346 4354
rect 15376 4676 15436 4715
rect 15376 4642 15389 4676
rect 15423 4642 15436 4676
rect 15376 4604 15436 4642
rect 15376 4570 15389 4604
rect 15423 4570 15436 4604
rect 15376 4532 15436 4570
rect 15376 4498 15389 4532
rect 15423 4498 15436 4532
rect 15376 4460 15436 4498
rect 15376 4426 15389 4460
rect 15423 4426 15436 4460
rect 15376 4388 15436 4426
rect 15376 4354 15389 4388
rect 15423 4354 15436 4388
rect 15376 4315 15436 4354
rect 15466 4676 15526 4715
rect 15466 4642 15479 4676
rect 15513 4642 15526 4676
rect 15466 4604 15526 4642
rect 15466 4570 15479 4604
rect 15513 4570 15526 4604
rect 15466 4532 15526 4570
rect 15466 4498 15479 4532
rect 15513 4498 15526 4532
rect 15466 4460 15526 4498
rect 15466 4426 15479 4460
rect 15513 4426 15526 4460
rect 15466 4388 15526 4426
rect 15466 4354 15479 4388
rect 15513 4354 15526 4388
rect 15466 4315 15526 4354
rect 15556 4676 15616 4715
rect 15556 4642 15569 4676
rect 15603 4642 15616 4676
rect 15556 4604 15616 4642
rect 15556 4570 15569 4604
rect 15603 4570 15616 4604
rect 15556 4532 15616 4570
rect 15556 4498 15569 4532
rect 15603 4498 15616 4532
rect 15556 4460 15616 4498
rect 15556 4426 15569 4460
rect 15603 4426 15616 4460
rect 15556 4388 15616 4426
rect 15556 4354 15569 4388
rect 15603 4354 15616 4388
rect 15556 4315 15616 4354
rect 24854 4676 24914 4715
rect 24854 4642 24867 4676
rect 24901 4642 24914 4676
rect 24854 4604 24914 4642
rect 24854 4570 24867 4604
rect 24901 4570 24914 4604
rect 24854 4532 24914 4570
rect 24854 4498 24867 4532
rect 24901 4498 24914 4532
rect 24854 4460 24914 4498
rect 24854 4426 24867 4460
rect 24901 4426 24914 4460
rect 24854 4388 24914 4426
rect 24854 4354 24867 4388
rect 24901 4354 24914 4388
rect 24854 4315 24914 4354
rect 24984 4676 25044 4715
rect 24984 4642 24997 4676
rect 25031 4642 25044 4676
rect 24984 4604 25044 4642
rect 24984 4570 24997 4604
rect 25031 4570 25044 4604
rect 24984 4532 25044 4570
rect 24984 4498 24997 4532
rect 25031 4498 25044 4532
rect 24984 4460 25044 4498
rect 24984 4426 24997 4460
rect 25031 4426 25044 4460
rect 24984 4388 25044 4426
rect 24984 4354 24997 4388
rect 25031 4354 25044 4388
rect 24984 4315 25044 4354
rect 25244 4676 25304 4715
rect 25244 4642 25257 4676
rect 25291 4642 25304 4676
rect 25244 4604 25304 4642
rect 25244 4570 25257 4604
rect 25291 4570 25304 4604
rect 25244 4532 25304 4570
rect 25244 4498 25257 4532
rect 25291 4498 25304 4532
rect 25244 4460 25304 4498
rect 25244 4426 25257 4460
rect 25291 4426 25304 4460
rect 25244 4388 25304 4426
rect 25244 4354 25257 4388
rect 25291 4354 25304 4388
rect 25244 4315 25304 4354
rect 25374 4676 25434 4715
rect 25374 4642 25387 4676
rect 25421 4642 25434 4676
rect 25374 4604 25434 4642
rect 25374 4570 25387 4604
rect 25421 4570 25434 4604
rect 25374 4532 25434 4570
rect 25374 4498 25387 4532
rect 25421 4498 25434 4532
rect 25374 4460 25434 4498
rect 25374 4426 25387 4460
rect 25421 4426 25434 4460
rect 25374 4388 25434 4426
rect 25374 4354 25387 4388
rect 25421 4354 25434 4388
rect 25374 4315 25434 4354
rect 25634 4676 25694 4715
rect 25634 4642 25647 4676
rect 25681 4642 25694 4676
rect 25634 4604 25694 4642
rect 25634 4570 25647 4604
rect 25681 4570 25694 4604
rect 25634 4532 25694 4570
rect 25634 4498 25647 4532
rect 25681 4498 25694 4532
rect 25634 4460 25694 4498
rect 25634 4426 25647 4460
rect 25681 4426 25694 4460
rect 25634 4388 25694 4426
rect 25634 4354 25647 4388
rect 25681 4354 25694 4388
rect 25634 4315 25694 4354
rect 25764 4676 25824 4715
rect 25764 4642 25777 4676
rect 25811 4642 25824 4676
rect 25764 4604 25824 4642
rect 25764 4570 25777 4604
rect 25811 4570 25824 4604
rect 25764 4532 25824 4570
rect 25764 4498 25777 4532
rect 25811 4498 25824 4532
rect 25764 4460 25824 4498
rect 25764 4426 25777 4460
rect 25811 4426 25824 4460
rect 25764 4388 25824 4426
rect 25764 4354 25777 4388
rect 25811 4354 25824 4388
rect 25764 4315 25824 4354
rect 26024 4676 26084 4715
rect 26024 4642 26037 4676
rect 26071 4642 26084 4676
rect 26024 4604 26084 4642
rect 26024 4570 26037 4604
rect 26071 4570 26084 4604
rect 26024 4532 26084 4570
rect 26024 4498 26037 4532
rect 26071 4498 26084 4532
rect 26024 4460 26084 4498
rect 26024 4426 26037 4460
rect 26071 4426 26084 4460
rect 26024 4388 26084 4426
rect 26024 4354 26037 4388
rect 26071 4354 26084 4388
rect 26024 4315 26084 4354
rect 26154 4676 26214 4715
rect 26154 4642 26167 4676
rect 26201 4642 26214 4676
rect 26154 4604 26214 4642
rect 26154 4570 26167 4604
rect 26201 4570 26214 4604
rect 26154 4532 26214 4570
rect 26154 4498 26167 4532
rect 26201 4498 26214 4532
rect 26154 4460 26214 4498
rect 26154 4426 26167 4460
rect 26201 4426 26214 4460
rect 26154 4388 26214 4426
rect 26154 4354 26167 4388
rect 26201 4354 26214 4388
rect 26154 4315 26214 4354
rect 26414 4676 26474 4715
rect 26414 4642 26427 4676
rect 26461 4642 26474 4676
rect 26414 4604 26474 4642
rect 26414 4570 26427 4604
rect 26461 4570 26474 4604
rect 26414 4532 26474 4570
rect 26414 4498 26427 4532
rect 26461 4498 26474 4532
rect 26414 4460 26474 4498
rect 26414 4426 26427 4460
rect 26461 4426 26474 4460
rect 26414 4388 26474 4426
rect 26414 4354 26427 4388
rect 26461 4354 26474 4388
rect 26414 4315 26474 4354
rect 26544 4676 26604 4715
rect 26544 4642 26557 4676
rect 26591 4642 26604 4676
rect 26544 4604 26604 4642
rect 26544 4570 26557 4604
rect 26591 4570 26604 4604
rect 26544 4532 26604 4570
rect 26544 4498 26557 4532
rect 26591 4498 26604 4532
rect 26544 4460 26604 4498
rect 26544 4426 26557 4460
rect 26591 4426 26604 4460
rect 26544 4388 26604 4426
rect 26544 4354 26557 4388
rect 26591 4354 26604 4388
rect 26544 4315 26604 4354
rect 26788 4676 26848 4715
rect 26788 4642 26801 4676
rect 26835 4642 26848 4676
rect 26788 4604 26848 4642
rect 26788 4570 26801 4604
rect 26835 4570 26848 4604
rect 26788 4532 26848 4570
rect 26788 4498 26801 4532
rect 26835 4498 26848 4532
rect 26788 4460 26848 4498
rect 26788 4426 26801 4460
rect 26835 4426 26848 4460
rect 26788 4388 26848 4426
rect 26788 4354 26801 4388
rect 26835 4354 26848 4388
rect 26788 4315 26848 4354
rect 26878 4676 26938 4715
rect 26878 4642 26891 4676
rect 26925 4642 26938 4676
rect 26878 4604 26938 4642
rect 26878 4570 26891 4604
rect 26925 4570 26938 4604
rect 26878 4532 26938 4570
rect 26878 4498 26891 4532
rect 26925 4498 26938 4532
rect 26878 4460 26938 4498
rect 26878 4426 26891 4460
rect 26925 4426 26938 4460
rect 26878 4388 26938 4426
rect 26878 4354 26891 4388
rect 26925 4354 26938 4388
rect 26878 4315 26938 4354
rect 26968 4676 27028 4715
rect 26968 4642 26981 4676
rect 27015 4642 27028 4676
rect 26968 4604 27028 4642
rect 26968 4570 26981 4604
rect 27015 4570 27028 4604
rect 26968 4532 27028 4570
rect 26968 4498 26981 4532
rect 27015 4498 27028 4532
rect 26968 4460 27028 4498
rect 26968 4426 26981 4460
rect 27015 4426 27028 4460
rect 26968 4388 27028 4426
rect 26968 4354 26981 4388
rect 27015 4354 27028 4388
rect 26968 4315 27028 4354
rect 27058 4676 27118 4715
rect 27058 4642 27071 4676
rect 27105 4642 27118 4676
rect 27058 4604 27118 4642
rect 27058 4570 27071 4604
rect 27105 4570 27118 4604
rect 27058 4532 27118 4570
rect 27058 4498 27071 4532
rect 27105 4498 27118 4532
rect 27058 4460 27118 4498
rect 27058 4426 27071 4460
rect 27105 4426 27118 4460
rect 27058 4388 27118 4426
rect 27058 4354 27071 4388
rect 27105 4354 27118 4388
rect 27058 4315 27118 4354
rect 27148 4676 27208 4715
rect 27148 4642 27161 4676
rect 27195 4642 27208 4676
rect 27148 4604 27208 4642
rect 27148 4570 27161 4604
rect 27195 4570 27208 4604
rect 27148 4532 27208 4570
rect 27148 4498 27161 4532
rect 27195 4498 27208 4532
rect 27148 4460 27208 4498
rect 27148 4426 27161 4460
rect 27195 4426 27208 4460
rect 27148 4388 27208 4426
rect 27148 4354 27161 4388
rect 27195 4354 27208 4388
rect 27148 4315 27208 4354
rect 13262 1872 13322 1911
rect 13262 1838 13275 1872
rect 13309 1838 13322 1872
rect 13262 1800 13322 1838
rect 13262 1766 13275 1800
rect 13309 1766 13322 1800
rect 13262 1728 13322 1766
rect 13262 1694 13275 1728
rect 13309 1694 13322 1728
rect 13262 1656 13322 1694
rect 13262 1622 13275 1656
rect 13309 1622 13322 1656
rect 13262 1584 13322 1622
rect 13262 1550 13275 1584
rect 13309 1550 13322 1584
rect 13262 1511 13322 1550
rect 13392 1872 13452 1911
rect 13392 1838 13405 1872
rect 13439 1838 13452 1872
rect 13392 1800 13452 1838
rect 13392 1766 13405 1800
rect 13439 1766 13452 1800
rect 13392 1728 13452 1766
rect 13392 1694 13405 1728
rect 13439 1694 13452 1728
rect 13392 1656 13452 1694
rect 13392 1622 13405 1656
rect 13439 1622 13452 1656
rect 13392 1584 13452 1622
rect 13392 1550 13405 1584
rect 13439 1550 13452 1584
rect 13392 1511 13452 1550
rect 13652 1872 13712 1911
rect 13652 1838 13665 1872
rect 13699 1838 13712 1872
rect 13652 1800 13712 1838
rect 13652 1766 13665 1800
rect 13699 1766 13712 1800
rect 13652 1728 13712 1766
rect 13652 1694 13665 1728
rect 13699 1694 13712 1728
rect 13652 1656 13712 1694
rect 13652 1622 13665 1656
rect 13699 1622 13712 1656
rect 13652 1584 13712 1622
rect 13652 1550 13665 1584
rect 13699 1550 13712 1584
rect 13652 1511 13712 1550
rect 13782 1872 13842 1911
rect 13782 1838 13795 1872
rect 13829 1838 13842 1872
rect 13782 1800 13842 1838
rect 13782 1766 13795 1800
rect 13829 1766 13842 1800
rect 13782 1728 13842 1766
rect 13782 1694 13795 1728
rect 13829 1694 13842 1728
rect 13782 1656 13842 1694
rect 13782 1622 13795 1656
rect 13829 1622 13842 1656
rect 13782 1584 13842 1622
rect 13782 1550 13795 1584
rect 13829 1550 13842 1584
rect 13782 1511 13842 1550
rect 14042 1872 14102 1911
rect 14042 1838 14055 1872
rect 14089 1838 14102 1872
rect 14042 1800 14102 1838
rect 14042 1766 14055 1800
rect 14089 1766 14102 1800
rect 14042 1728 14102 1766
rect 14042 1694 14055 1728
rect 14089 1694 14102 1728
rect 14042 1656 14102 1694
rect 14042 1622 14055 1656
rect 14089 1622 14102 1656
rect 14042 1584 14102 1622
rect 14042 1550 14055 1584
rect 14089 1550 14102 1584
rect 14042 1511 14102 1550
rect 14172 1872 14232 1911
rect 14172 1838 14185 1872
rect 14219 1838 14232 1872
rect 14172 1800 14232 1838
rect 14172 1766 14185 1800
rect 14219 1766 14232 1800
rect 14172 1728 14232 1766
rect 14172 1694 14185 1728
rect 14219 1694 14232 1728
rect 14172 1656 14232 1694
rect 14172 1622 14185 1656
rect 14219 1622 14232 1656
rect 14172 1584 14232 1622
rect 14172 1550 14185 1584
rect 14219 1550 14232 1584
rect 14172 1511 14232 1550
rect 14432 1872 14492 1911
rect 14432 1838 14445 1872
rect 14479 1838 14492 1872
rect 14432 1800 14492 1838
rect 14432 1766 14445 1800
rect 14479 1766 14492 1800
rect 14432 1728 14492 1766
rect 14432 1694 14445 1728
rect 14479 1694 14492 1728
rect 14432 1656 14492 1694
rect 14432 1622 14445 1656
rect 14479 1622 14492 1656
rect 14432 1584 14492 1622
rect 14432 1550 14445 1584
rect 14479 1550 14492 1584
rect 14432 1511 14492 1550
rect 14562 1872 14622 1911
rect 14562 1838 14575 1872
rect 14609 1838 14622 1872
rect 14562 1800 14622 1838
rect 14562 1766 14575 1800
rect 14609 1766 14622 1800
rect 14562 1728 14622 1766
rect 14562 1694 14575 1728
rect 14609 1694 14622 1728
rect 14562 1656 14622 1694
rect 14562 1622 14575 1656
rect 14609 1622 14622 1656
rect 14562 1584 14622 1622
rect 14562 1550 14575 1584
rect 14609 1550 14622 1584
rect 14562 1511 14622 1550
rect 14822 1872 14882 1911
rect 14822 1838 14835 1872
rect 14869 1838 14882 1872
rect 14822 1800 14882 1838
rect 14822 1766 14835 1800
rect 14869 1766 14882 1800
rect 14822 1728 14882 1766
rect 14822 1694 14835 1728
rect 14869 1694 14882 1728
rect 14822 1656 14882 1694
rect 14822 1622 14835 1656
rect 14869 1622 14882 1656
rect 14822 1584 14882 1622
rect 14822 1550 14835 1584
rect 14869 1550 14882 1584
rect 14822 1511 14882 1550
rect 14952 1872 15012 1911
rect 14952 1838 14965 1872
rect 14999 1838 15012 1872
rect 14952 1800 15012 1838
rect 14952 1766 14965 1800
rect 14999 1766 15012 1800
rect 14952 1728 15012 1766
rect 14952 1694 14965 1728
rect 14999 1694 15012 1728
rect 14952 1656 15012 1694
rect 14952 1622 14965 1656
rect 14999 1622 15012 1656
rect 14952 1584 15012 1622
rect 14952 1550 14965 1584
rect 14999 1550 15012 1584
rect 14952 1511 15012 1550
rect 15212 1872 15272 1911
rect 15212 1838 15225 1872
rect 15259 1838 15272 1872
rect 15212 1800 15272 1838
rect 15212 1766 15225 1800
rect 15259 1766 15272 1800
rect 15212 1728 15272 1766
rect 15212 1694 15225 1728
rect 15259 1694 15272 1728
rect 15212 1656 15272 1694
rect 15212 1622 15225 1656
rect 15259 1622 15272 1656
rect 15212 1584 15272 1622
rect 15212 1550 15225 1584
rect 15259 1550 15272 1584
rect 15212 1511 15272 1550
rect 15342 1872 15402 1911
rect 15342 1838 15355 1872
rect 15389 1838 15402 1872
rect 15342 1800 15402 1838
rect 15342 1766 15355 1800
rect 15389 1766 15402 1800
rect 15342 1728 15402 1766
rect 15342 1694 15355 1728
rect 15389 1694 15402 1728
rect 15342 1656 15402 1694
rect 15342 1622 15355 1656
rect 15389 1622 15402 1656
rect 15342 1584 15402 1622
rect 15342 1550 15355 1584
rect 15389 1550 15402 1584
rect 15342 1511 15402 1550
rect 24854 1872 24914 1911
rect 24854 1838 24867 1872
rect 24901 1838 24914 1872
rect 24854 1800 24914 1838
rect 24854 1766 24867 1800
rect 24901 1766 24914 1800
rect 24854 1728 24914 1766
rect 24854 1694 24867 1728
rect 24901 1694 24914 1728
rect 24854 1656 24914 1694
rect 24854 1622 24867 1656
rect 24901 1622 24914 1656
rect 24854 1584 24914 1622
rect 24854 1550 24867 1584
rect 24901 1550 24914 1584
rect 24854 1511 24914 1550
rect 24984 1872 25044 1911
rect 24984 1838 24997 1872
rect 25031 1838 25044 1872
rect 24984 1800 25044 1838
rect 24984 1766 24997 1800
rect 25031 1766 25044 1800
rect 24984 1728 25044 1766
rect 24984 1694 24997 1728
rect 25031 1694 25044 1728
rect 24984 1656 25044 1694
rect 24984 1622 24997 1656
rect 25031 1622 25044 1656
rect 24984 1584 25044 1622
rect 24984 1550 24997 1584
rect 25031 1550 25044 1584
rect 24984 1511 25044 1550
rect 25244 1872 25304 1911
rect 25244 1838 25257 1872
rect 25291 1838 25304 1872
rect 25244 1800 25304 1838
rect 25244 1766 25257 1800
rect 25291 1766 25304 1800
rect 25244 1728 25304 1766
rect 25244 1694 25257 1728
rect 25291 1694 25304 1728
rect 25244 1656 25304 1694
rect 25244 1622 25257 1656
rect 25291 1622 25304 1656
rect 25244 1584 25304 1622
rect 25244 1550 25257 1584
rect 25291 1550 25304 1584
rect 25244 1511 25304 1550
rect 25374 1872 25434 1911
rect 25374 1838 25387 1872
rect 25421 1838 25434 1872
rect 25374 1800 25434 1838
rect 25374 1766 25387 1800
rect 25421 1766 25434 1800
rect 25374 1728 25434 1766
rect 25374 1694 25387 1728
rect 25421 1694 25434 1728
rect 25374 1656 25434 1694
rect 25374 1622 25387 1656
rect 25421 1622 25434 1656
rect 25374 1584 25434 1622
rect 25374 1550 25387 1584
rect 25421 1550 25434 1584
rect 25374 1511 25434 1550
rect 25634 1872 25694 1911
rect 25634 1838 25647 1872
rect 25681 1838 25694 1872
rect 25634 1800 25694 1838
rect 25634 1766 25647 1800
rect 25681 1766 25694 1800
rect 25634 1728 25694 1766
rect 25634 1694 25647 1728
rect 25681 1694 25694 1728
rect 25634 1656 25694 1694
rect 25634 1622 25647 1656
rect 25681 1622 25694 1656
rect 25634 1584 25694 1622
rect 25634 1550 25647 1584
rect 25681 1550 25694 1584
rect 25634 1511 25694 1550
rect 25764 1872 25824 1911
rect 25764 1838 25777 1872
rect 25811 1838 25824 1872
rect 25764 1800 25824 1838
rect 25764 1766 25777 1800
rect 25811 1766 25824 1800
rect 25764 1728 25824 1766
rect 25764 1694 25777 1728
rect 25811 1694 25824 1728
rect 25764 1656 25824 1694
rect 25764 1622 25777 1656
rect 25811 1622 25824 1656
rect 25764 1584 25824 1622
rect 25764 1550 25777 1584
rect 25811 1550 25824 1584
rect 25764 1511 25824 1550
rect 26024 1872 26084 1911
rect 26024 1838 26037 1872
rect 26071 1838 26084 1872
rect 26024 1800 26084 1838
rect 26024 1766 26037 1800
rect 26071 1766 26084 1800
rect 26024 1728 26084 1766
rect 26024 1694 26037 1728
rect 26071 1694 26084 1728
rect 26024 1656 26084 1694
rect 26024 1622 26037 1656
rect 26071 1622 26084 1656
rect 26024 1584 26084 1622
rect 26024 1550 26037 1584
rect 26071 1550 26084 1584
rect 26024 1511 26084 1550
rect 26154 1872 26214 1911
rect 26154 1838 26167 1872
rect 26201 1838 26214 1872
rect 26154 1800 26214 1838
rect 26154 1766 26167 1800
rect 26201 1766 26214 1800
rect 26154 1728 26214 1766
rect 26154 1694 26167 1728
rect 26201 1694 26214 1728
rect 26154 1656 26214 1694
rect 26154 1622 26167 1656
rect 26201 1622 26214 1656
rect 26154 1584 26214 1622
rect 26154 1550 26167 1584
rect 26201 1550 26214 1584
rect 26154 1511 26214 1550
rect 26414 1872 26474 1911
rect 26414 1838 26427 1872
rect 26461 1838 26474 1872
rect 26414 1800 26474 1838
rect 26414 1766 26427 1800
rect 26461 1766 26474 1800
rect 26414 1728 26474 1766
rect 26414 1694 26427 1728
rect 26461 1694 26474 1728
rect 26414 1656 26474 1694
rect 26414 1622 26427 1656
rect 26461 1622 26474 1656
rect 26414 1584 26474 1622
rect 26414 1550 26427 1584
rect 26461 1550 26474 1584
rect 26414 1511 26474 1550
rect 26544 1872 26604 1911
rect 26544 1838 26557 1872
rect 26591 1838 26604 1872
rect 26544 1800 26604 1838
rect 26544 1766 26557 1800
rect 26591 1766 26604 1800
rect 26544 1728 26604 1766
rect 26544 1694 26557 1728
rect 26591 1694 26604 1728
rect 26544 1656 26604 1694
rect 26544 1622 26557 1656
rect 26591 1622 26604 1656
rect 26544 1584 26604 1622
rect 26544 1550 26557 1584
rect 26591 1550 26604 1584
rect 26544 1511 26604 1550
rect 26804 1872 26864 1911
rect 26804 1838 26817 1872
rect 26851 1838 26864 1872
rect 26804 1800 26864 1838
rect 26804 1766 26817 1800
rect 26851 1766 26864 1800
rect 26804 1728 26864 1766
rect 26804 1694 26817 1728
rect 26851 1694 26864 1728
rect 26804 1656 26864 1694
rect 26804 1622 26817 1656
rect 26851 1622 26864 1656
rect 26804 1584 26864 1622
rect 26804 1550 26817 1584
rect 26851 1550 26864 1584
rect 26804 1511 26864 1550
rect 26934 1872 26994 1911
rect 26934 1838 26947 1872
rect 26981 1838 26994 1872
rect 26934 1800 26994 1838
rect 26934 1766 26947 1800
rect 26981 1766 26994 1800
rect 26934 1728 26994 1766
rect 26934 1694 26947 1728
rect 26981 1694 26994 1728
rect 26934 1656 26994 1694
rect 26934 1622 26947 1656
rect 26981 1622 26994 1656
rect 26934 1584 26994 1622
rect 26934 1550 26947 1584
rect 26981 1550 26994 1584
rect 26934 1511 26994 1550
rect 13132 1324 13192 1363
rect 13132 1290 13145 1324
rect 13179 1290 13192 1324
rect 13132 1252 13192 1290
rect 13132 1218 13145 1252
rect 13179 1218 13192 1252
rect 13132 1180 13192 1218
rect 13132 1146 13145 1180
rect 13179 1146 13192 1180
rect 13132 1108 13192 1146
rect 13132 1074 13145 1108
rect 13179 1074 13192 1108
rect 13132 1036 13192 1074
rect 13132 1002 13145 1036
rect 13179 1002 13192 1036
rect 13132 963 13192 1002
rect 13262 1324 13322 1363
rect 13262 1290 13275 1324
rect 13309 1290 13322 1324
rect 13262 1252 13322 1290
rect 13262 1218 13275 1252
rect 13309 1218 13322 1252
rect 13262 1180 13322 1218
rect 13262 1146 13275 1180
rect 13309 1146 13322 1180
rect 13262 1108 13322 1146
rect 13262 1074 13275 1108
rect 13309 1074 13322 1108
rect 13262 1036 13322 1074
rect 13262 1002 13275 1036
rect 13309 1002 13322 1036
rect 13262 963 13322 1002
rect 13392 1324 13452 1363
rect 13392 1290 13405 1324
rect 13439 1290 13452 1324
rect 13392 1252 13452 1290
rect 13392 1218 13405 1252
rect 13439 1218 13452 1252
rect 13392 1180 13452 1218
rect 13392 1146 13405 1180
rect 13439 1146 13452 1180
rect 13392 1108 13452 1146
rect 13392 1074 13405 1108
rect 13439 1074 13452 1108
rect 13392 1036 13452 1074
rect 13392 1002 13405 1036
rect 13439 1002 13452 1036
rect 13392 963 13452 1002
rect 13522 1324 13582 1363
rect 13522 1290 13535 1324
rect 13569 1290 13582 1324
rect 13522 1252 13582 1290
rect 13522 1218 13535 1252
rect 13569 1218 13582 1252
rect 13522 1180 13582 1218
rect 13522 1146 13535 1180
rect 13569 1146 13582 1180
rect 13522 1108 13582 1146
rect 13522 1074 13535 1108
rect 13569 1074 13582 1108
rect 13522 1036 13582 1074
rect 13522 1002 13535 1036
rect 13569 1002 13582 1036
rect 13522 963 13582 1002
rect 13652 1324 13712 1363
rect 13652 1290 13665 1324
rect 13699 1290 13712 1324
rect 13652 1252 13712 1290
rect 13652 1218 13665 1252
rect 13699 1218 13712 1252
rect 13652 1180 13712 1218
rect 13652 1146 13665 1180
rect 13699 1146 13712 1180
rect 13652 1108 13712 1146
rect 13652 1074 13665 1108
rect 13699 1074 13712 1108
rect 13652 1036 13712 1074
rect 13652 1002 13665 1036
rect 13699 1002 13712 1036
rect 13652 963 13712 1002
rect 13782 1324 13842 1363
rect 13782 1290 13795 1324
rect 13829 1290 13842 1324
rect 13782 1252 13842 1290
rect 13782 1218 13795 1252
rect 13829 1218 13842 1252
rect 13782 1180 13842 1218
rect 13782 1146 13795 1180
rect 13829 1146 13842 1180
rect 13782 1108 13842 1146
rect 13782 1074 13795 1108
rect 13829 1074 13842 1108
rect 13782 1036 13842 1074
rect 13782 1002 13795 1036
rect 13829 1002 13842 1036
rect 13782 963 13842 1002
rect 13912 1324 13972 1363
rect 13912 1290 13925 1324
rect 13959 1290 13972 1324
rect 13912 1252 13972 1290
rect 13912 1218 13925 1252
rect 13959 1218 13972 1252
rect 13912 1180 13972 1218
rect 13912 1146 13925 1180
rect 13959 1146 13972 1180
rect 13912 1108 13972 1146
rect 13912 1074 13925 1108
rect 13959 1074 13972 1108
rect 13912 1036 13972 1074
rect 13912 1002 13925 1036
rect 13959 1002 13972 1036
rect 13912 963 13972 1002
rect 14042 1324 14102 1363
rect 14042 1290 14055 1324
rect 14089 1290 14102 1324
rect 14042 1252 14102 1290
rect 14042 1218 14055 1252
rect 14089 1218 14102 1252
rect 14042 1180 14102 1218
rect 14042 1146 14055 1180
rect 14089 1146 14102 1180
rect 14042 1108 14102 1146
rect 14042 1074 14055 1108
rect 14089 1074 14102 1108
rect 14042 1036 14102 1074
rect 14042 1002 14055 1036
rect 14089 1002 14102 1036
rect 14042 963 14102 1002
rect 14172 1324 14232 1363
rect 14172 1290 14185 1324
rect 14219 1290 14232 1324
rect 14172 1252 14232 1290
rect 14172 1218 14185 1252
rect 14219 1218 14232 1252
rect 14172 1180 14232 1218
rect 14172 1146 14185 1180
rect 14219 1146 14232 1180
rect 14172 1108 14232 1146
rect 14172 1074 14185 1108
rect 14219 1074 14232 1108
rect 14172 1036 14232 1074
rect 14172 1002 14185 1036
rect 14219 1002 14232 1036
rect 14172 963 14232 1002
rect 14302 1324 14362 1363
rect 14302 1290 14315 1324
rect 14349 1290 14362 1324
rect 14302 1252 14362 1290
rect 14302 1218 14315 1252
rect 14349 1218 14362 1252
rect 14302 1180 14362 1218
rect 14302 1146 14315 1180
rect 14349 1146 14362 1180
rect 14302 1108 14362 1146
rect 14302 1074 14315 1108
rect 14349 1074 14362 1108
rect 14302 1036 14362 1074
rect 14302 1002 14315 1036
rect 14349 1002 14362 1036
rect 14302 963 14362 1002
rect 14432 1324 14492 1363
rect 14432 1290 14445 1324
rect 14479 1290 14492 1324
rect 14432 1252 14492 1290
rect 14432 1218 14445 1252
rect 14479 1218 14492 1252
rect 14432 1180 14492 1218
rect 14432 1146 14445 1180
rect 14479 1146 14492 1180
rect 14432 1108 14492 1146
rect 14432 1074 14445 1108
rect 14479 1074 14492 1108
rect 14432 1036 14492 1074
rect 14432 1002 14445 1036
rect 14479 1002 14492 1036
rect 14432 963 14492 1002
rect 14562 1324 14622 1363
rect 14562 1290 14575 1324
rect 14609 1290 14622 1324
rect 14562 1252 14622 1290
rect 14562 1218 14575 1252
rect 14609 1218 14622 1252
rect 14562 1180 14622 1218
rect 14562 1146 14575 1180
rect 14609 1146 14622 1180
rect 14562 1108 14622 1146
rect 14562 1074 14575 1108
rect 14609 1074 14622 1108
rect 14562 1036 14622 1074
rect 14562 1002 14575 1036
rect 14609 1002 14622 1036
rect 14562 963 14622 1002
rect 14692 1324 14752 1363
rect 14692 1290 14705 1324
rect 14739 1290 14752 1324
rect 14692 1252 14752 1290
rect 14692 1218 14705 1252
rect 14739 1218 14752 1252
rect 14692 1180 14752 1218
rect 14692 1146 14705 1180
rect 14739 1146 14752 1180
rect 14692 1108 14752 1146
rect 14692 1074 14705 1108
rect 14739 1074 14752 1108
rect 14692 1036 14752 1074
rect 14692 1002 14705 1036
rect 14739 1002 14752 1036
rect 14692 963 14752 1002
rect 14822 1324 14882 1363
rect 14822 1290 14835 1324
rect 14869 1290 14882 1324
rect 14822 1252 14882 1290
rect 14822 1218 14835 1252
rect 14869 1218 14882 1252
rect 14822 1180 14882 1218
rect 14822 1146 14835 1180
rect 14869 1146 14882 1180
rect 14822 1108 14882 1146
rect 14822 1074 14835 1108
rect 14869 1074 14882 1108
rect 14822 1036 14882 1074
rect 14822 1002 14835 1036
rect 14869 1002 14882 1036
rect 14822 963 14882 1002
rect 14952 1324 15012 1363
rect 14952 1290 14965 1324
rect 14999 1290 15012 1324
rect 14952 1252 15012 1290
rect 14952 1218 14965 1252
rect 14999 1218 15012 1252
rect 14952 1180 15012 1218
rect 14952 1146 14965 1180
rect 14999 1146 15012 1180
rect 14952 1108 15012 1146
rect 14952 1074 14965 1108
rect 14999 1074 15012 1108
rect 14952 1036 15012 1074
rect 14952 1002 14965 1036
rect 14999 1002 15012 1036
rect 14952 963 15012 1002
rect 15082 1324 15142 1363
rect 15082 1290 15095 1324
rect 15129 1290 15142 1324
rect 15082 1252 15142 1290
rect 15082 1218 15095 1252
rect 15129 1218 15142 1252
rect 15082 1180 15142 1218
rect 15082 1146 15095 1180
rect 15129 1146 15142 1180
rect 15082 1108 15142 1146
rect 15082 1074 15095 1108
rect 15129 1074 15142 1108
rect 15082 1036 15142 1074
rect 15082 1002 15095 1036
rect 15129 1002 15142 1036
rect 15082 963 15142 1002
rect 15212 1324 15272 1363
rect 15212 1290 15225 1324
rect 15259 1290 15272 1324
rect 15212 1252 15272 1290
rect 15212 1218 15225 1252
rect 15259 1218 15272 1252
rect 15212 1180 15272 1218
rect 15212 1146 15225 1180
rect 15259 1146 15272 1180
rect 15212 1108 15272 1146
rect 15212 1074 15225 1108
rect 15259 1074 15272 1108
rect 15212 1036 15272 1074
rect 15212 1002 15225 1036
rect 15259 1002 15272 1036
rect 15212 963 15272 1002
rect 15342 1324 15402 1363
rect 15342 1290 15355 1324
rect 15389 1290 15402 1324
rect 15342 1252 15402 1290
rect 15342 1218 15355 1252
rect 15389 1218 15402 1252
rect 15342 1180 15402 1218
rect 15342 1146 15355 1180
rect 15389 1146 15402 1180
rect 15342 1108 15402 1146
rect 15342 1074 15355 1108
rect 15389 1074 15402 1108
rect 15342 1036 15402 1074
rect 15342 1002 15355 1036
rect 15389 1002 15402 1036
rect 15342 963 15402 1002
rect 15472 1324 15532 1363
rect 15472 1290 15485 1324
rect 15519 1290 15532 1324
rect 15472 1252 15532 1290
rect 15472 1218 15485 1252
rect 15519 1218 15532 1252
rect 15472 1180 15532 1218
rect 15472 1146 15485 1180
rect 15519 1146 15532 1180
rect 15472 1108 15532 1146
rect 15472 1074 15485 1108
rect 15519 1074 15532 1108
rect 15472 1036 15532 1074
rect 15472 1002 15485 1036
rect 15519 1002 15532 1036
rect 15472 963 15532 1002
rect 24724 1324 24784 1363
rect 24724 1290 24737 1324
rect 24771 1290 24784 1324
rect 24724 1252 24784 1290
rect 24724 1218 24737 1252
rect 24771 1218 24784 1252
rect 24724 1180 24784 1218
rect 24724 1146 24737 1180
rect 24771 1146 24784 1180
rect 24724 1108 24784 1146
rect 24724 1074 24737 1108
rect 24771 1074 24784 1108
rect 24724 1036 24784 1074
rect 24724 1002 24737 1036
rect 24771 1002 24784 1036
rect 24724 963 24784 1002
rect 24854 1324 24914 1363
rect 24854 1290 24867 1324
rect 24901 1290 24914 1324
rect 24854 1252 24914 1290
rect 24854 1218 24867 1252
rect 24901 1218 24914 1252
rect 24854 1180 24914 1218
rect 24854 1146 24867 1180
rect 24901 1146 24914 1180
rect 24854 1108 24914 1146
rect 24854 1074 24867 1108
rect 24901 1074 24914 1108
rect 24854 1036 24914 1074
rect 24854 1002 24867 1036
rect 24901 1002 24914 1036
rect 24854 963 24914 1002
rect 24984 1324 25044 1363
rect 24984 1290 24997 1324
rect 25031 1290 25044 1324
rect 24984 1252 25044 1290
rect 24984 1218 24997 1252
rect 25031 1218 25044 1252
rect 24984 1180 25044 1218
rect 24984 1146 24997 1180
rect 25031 1146 25044 1180
rect 24984 1108 25044 1146
rect 24984 1074 24997 1108
rect 25031 1074 25044 1108
rect 24984 1036 25044 1074
rect 24984 1002 24997 1036
rect 25031 1002 25044 1036
rect 24984 963 25044 1002
rect 25114 1324 25174 1363
rect 25114 1290 25127 1324
rect 25161 1290 25174 1324
rect 25114 1252 25174 1290
rect 25114 1218 25127 1252
rect 25161 1218 25174 1252
rect 25114 1180 25174 1218
rect 25114 1146 25127 1180
rect 25161 1146 25174 1180
rect 25114 1108 25174 1146
rect 25114 1074 25127 1108
rect 25161 1074 25174 1108
rect 25114 1036 25174 1074
rect 25114 1002 25127 1036
rect 25161 1002 25174 1036
rect 25114 963 25174 1002
rect 25244 1324 25304 1363
rect 25244 1290 25257 1324
rect 25291 1290 25304 1324
rect 25244 1252 25304 1290
rect 25244 1218 25257 1252
rect 25291 1218 25304 1252
rect 25244 1180 25304 1218
rect 25244 1146 25257 1180
rect 25291 1146 25304 1180
rect 25244 1108 25304 1146
rect 25244 1074 25257 1108
rect 25291 1074 25304 1108
rect 25244 1036 25304 1074
rect 25244 1002 25257 1036
rect 25291 1002 25304 1036
rect 25244 963 25304 1002
rect 25374 1324 25434 1363
rect 25374 1290 25387 1324
rect 25421 1290 25434 1324
rect 25374 1252 25434 1290
rect 25374 1218 25387 1252
rect 25421 1218 25434 1252
rect 25374 1180 25434 1218
rect 25374 1146 25387 1180
rect 25421 1146 25434 1180
rect 25374 1108 25434 1146
rect 25374 1074 25387 1108
rect 25421 1074 25434 1108
rect 25374 1036 25434 1074
rect 25374 1002 25387 1036
rect 25421 1002 25434 1036
rect 25374 963 25434 1002
rect 25504 1324 25564 1363
rect 25504 1290 25517 1324
rect 25551 1290 25564 1324
rect 25504 1252 25564 1290
rect 25504 1218 25517 1252
rect 25551 1218 25564 1252
rect 25504 1180 25564 1218
rect 25504 1146 25517 1180
rect 25551 1146 25564 1180
rect 25504 1108 25564 1146
rect 25504 1074 25517 1108
rect 25551 1074 25564 1108
rect 25504 1036 25564 1074
rect 25504 1002 25517 1036
rect 25551 1002 25564 1036
rect 25504 963 25564 1002
rect 25634 1324 25694 1363
rect 25634 1290 25647 1324
rect 25681 1290 25694 1324
rect 25634 1252 25694 1290
rect 25634 1218 25647 1252
rect 25681 1218 25694 1252
rect 25634 1180 25694 1218
rect 25634 1146 25647 1180
rect 25681 1146 25694 1180
rect 25634 1108 25694 1146
rect 25634 1074 25647 1108
rect 25681 1074 25694 1108
rect 25634 1036 25694 1074
rect 25634 1002 25647 1036
rect 25681 1002 25694 1036
rect 25634 963 25694 1002
rect 25764 1324 25824 1363
rect 25764 1290 25777 1324
rect 25811 1290 25824 1324
rect 25764 1252 25824 1290
rect 25764 1218 25777 1252
rect 25811 1218 25824 1252
rect 25764 1180 25824 1218
rect 25764 1146 25777 1180
rect 25811 1146 25824 1180
rect 25764 1108 25824 1146
rect 25764 1074 25777 1108
rect 25811 1074 25824 1108
rect 25764 1036 25824 1074
rect 25764 1002 25777 1036
rect 25811 1002 25824 1036
rect 25764 963 25824 1002
rect 25894 1324 25954 1363
rect 25894 1290 25907 1324
rect 25941 1290 25954 1324
rect 25894 1252 25954 1290
rect 25894 1218 25907 1252
rect 25941 1218 25954 1252
rect 25894 1180 25954 1218
rect 25894 1146 25907 1180
rect 25941 1146 25954 1180
rect 25894 1108 25954 1146
rect 25894 1074 25907 1108
rect 25941 1074 25954 1108
rect 25894 1036 25954 1074
rect 25894 1002 25907 1036
rect 25941 1002 25954 1036
rect 25894 963 25954 1002
rect 26024 1324 26084 1363
rect 26024 1290 26037 1324
rect 26071 1290 26084 1324
rect 26024 1252 26084 1290
rect 26024 1218 26037 1252
rect 26071 1218 26084 1252
rect 26024 1180 26084 1218
rect 26024 1146 26037 1180
rect 26071 1146 26084 1180
rect 26024 1108 26084 1146
rect 26024 1074 26037 1108
rect 26071 1074 26084 1108
rect 26024 1036 26084 1074
rect 26024 1002 26037 1036
rect 26071 1002 26084 1036
rect 26024 963 26084 1002
rect 26154 1324 26214 1363
rect 26154 1290 26167 1324
rect 26201 1290 26214 1324
rect 26154 1252 26214 1290
rect 26154 1218 26167 1252
rect 26201 1218 26214 1252
rect 26154 1180 26214 1218
rect 26154 1146 26167 1180
rect 26201 1146 26214 1180
rect 26154 1108 26214 1146
rect 26154 1074 26167 1108
rect 26201 1074 26214 1108
rect 26154 1036 26214 1074
rect 26154 1002 26167 1036
rect 26201 1002 26214 1036
rect 26154 963 26214 1002
rect 26284 1324 26344 1363
rect 26284 1290 26297 1324
rect 26331 1290 26344 1324
rect 26284 1252 26344 1290
rect 26284 1218 26297 1252
rect 26331 1218 26344 1252
rect 26284 1180 26344 1218
rect 26284 1146 26297 1180
rect 26331 1146 26344 1180
rect 26284 1108 26344 1146
rect 26284 1074 26297 1108
rect 26331 1074 26344 1108
rect 26284 1036 26344 1074
rect 26284 1002 26297 1036
rect 26331 1002 26344 1036
rect 26284 963 26344 1002
rect 26414 1324 26474 1363
rect 26414 1290 26427 1324
rect 26461 1290 26474 1324
rect 26414 1252 26474 1290
rect 26414 1218 26427 1252
rect 26461 1218 26474 1252
rect 26414 1180 26474 1218
rect 26414 1146 26427 1180
rect 26461 1146 26474 1180
rect 26414 1108 26474 1146
rect 26414 1074 26427 1108
rect 26461 1074 26474 1108
rect 26414 1036 26474 1074
rect 26414 1002 26427 1036
rect 26461 1002 26474 1036
rect 26414 963 26474 1002
rect 26544 1324 26604 1363
rect 26544 1290 26557 1324
rect 26591 1290 26604 1324
rect 26544 1252 26604 1290
rect 26544 1218 26557 1252
rect 26591 1218 26604 1252
rect 26544 1180 26604 1218
rect 26544 1146 26557 1180
rect 26591 1146 26604 1180
rect 26544 1108 26604 1146
rect 26544 1074 26557 1108
rect 26591 1074 26604 1108
rect 26544 1036 26604 1074
rect 26544 1002 26557 1036
rect 26591 1002 26604 1036
rect 26544 963 26604 1002
rect 26674 1324 26734 1363
rect 26674 1290 26687 1324
rect 26721 1290 26734 1324
rect 26674 1252 26734 1290
rect 26674 1218 26687 1252
rect 26721 1218 26734 1252
rect 26674 1180 26734 1218
rect 26674 1146 26687 1180
rect 26721 1146 26734 1180
rect 26674 1108 26734 1146
rect 26674 1074 26687 1108
rect 26721 1074 26734 1108
rect 26674 1036 26734 1074
rect 26674 1002 26687 1036
rect 26721 1002 26734 1036
rect 26674 963 26734 1002
rect 26804 1324 26864 1363
rect 26804 1290 26817 1324
rect 26851 1290 26864 1324
rect 26804 1252 26864 1290
rect 26804 1218 26817 1252
rect 26851 1218 26864 1252
rect 26804 1180 26864 1218
rect 26804 1146 26817 1180
rect 26851 1146 26864 1180
rect 26804 1108 26864 1146
rect 26804 1074 26817 1108
rect 26851 1074 26864 1108
rect 26804 1036 26864 1074
rect 26804 1002 26817 1036
rect 26851 1002 26864 1036
rect 26804 963 26864 1002
rect 26934 1324 26994 1363
rect 26934 1290 26947 1324
rect 26981 1290 26994 1324
rect 26934 1252 26994 1290
rect 26934 1218 26947 1252
rect 26981 1218 26994 1252
rect 26934 1180 26994 1218
rect 26934 1146 26947 1180
rect 26981 1146 26994 1180
rect 26934 1108 26994 1146
rect 26934 1074 26947 1108
rect 26981 1074 26994 1108
rect 26934 1036 26994 1074
rect 26934 1002 26947 1036
rect 26981 1002 26994 1036
rect 26934 963 26994 1002
rect 27064 1324 27124 1363
rect 27064 1290 27077 1324
rect 27111 1290 27124 1324
rect 27064 1252 27124 1290
rect 27064 1218 27077 1252
rect 27111 1218 27124 1252
rect 27064 1180 27124 1218
rect 27064 1146 27077 1180
rect 27111 1146 27124 1180
rect 27064 1108 27124 1146
rect 27064 1074 27077 1108
rect 27111 1074 27124 1108
rect 27064 1036 27124 1074
rect 27064 1002 27077 1036
rect 27111 1002 27124 1036
rect 27064 963 27124 1002
<< ndiffc >>
rect 13275 3786 13309 3820
rect 13275 3714 13309 3748
rect 13405 3786 13439 3820
rect 13405 3714 13439 3748
rect 13535 3786 13569 3820
rect 13535 3714 13569 3748
rect 13665 3786 13699 3820
rect 13665 3714 13699 3748
rect 13795 3786 13829 3820
rect 13795 3714 13829 3748
rect 13925 3786 13959 3820
rect 13925 3714 13959 3748
rect 14055 3786 14089 3820
rect 14055 3714 14089 3748
rect 14185 3786 14219 3820
rect 14185 3714 14219 3748
rect 14315 3786 14349 3820
rect 14315 3714 14349 3748
rect 14445 3786 14479 3820
rect 14445 3714 14479 3748
rect 14575 3786 14609 3820
rect 14575 3714 14609 3748
rect 14705 3786 14739 3820
rect 14705 3714 14739 3748
rect 14835 3786 14869 3820
rect 14835 3714 14869 3748
rect 14965 3786 14999 3820
rect 14965 3714 14999 3748
rect 15095 3786 15129 3820
rect 15095 3714 15129 3748
rect 15209 3786 15243 3820
rect 15209 3714 15243 3748
rect 15299 3786 15333 3820
rect 15299 3714 15333 3748
rect 15389 3786 15423 3820
rect 15389 3714 15423 3748
rect 15479 3786 15513 3820
rect 15479 3714 15513 3748
rect 15569 3786 15603 3820
rect 15569 3714 15603 3748
rect 24867 3786 24901 3820
rect 24867 3714 24901 3748
rect 24997 3786 25031 3820
rect 24997 3714 25031 3748
rect 25127 3786 25161 3820
rect 25127 3714 25161 3748
rect 25257 3786 25291 3820
rect 25257 3714 25291 3748
rect 25387 3786 25421 3820
rect 25387 3714 25421 3748
rect 25517 3786 25551 3820
rect 25517 3714 25551 3748
rect 25647 3786 25681 3820
rect 25647 3714 25681 3748
rect 25777 3786 25811 3820
rect 25777 3714 25811 3748
rect 25907 3786 25941 3820
rect 25907 3714 25941 3748
rect 26037 3786 26071 3820
rect 26037 3714 26071 3748
rect 26167 3786 26201 3820
rect 26167 3714 26201 3748
rect 26297 3786 26331 3820
rect 26297 3714 26331 3748
rect 26427 3786 26461 3820
rect 26427 3714 26461 3748
rect 26557 3786 26591 3820
rect 26557 3714 26591 3748
rect 26687 3786 26721 3820
rect 26687 3714 26721 3748
rect 26801 3786 26835 3820
rect 26801 3714 26835 3748
rect 26891 3786 26925 3820
rect 26891 3714 26925 3748
rect 26981 3786 27015 3820
rect 26981 3714 27015 3748
rect 27071 3786 27105 3820
rect 27071 3714 27105 3748
rect 27161 3786 27195 3820
rect 27161 3714 27195 3748
rect 13015 3438 13049 3472
rect 13015 3366 13049 3400
rect 13145 3438 13179 3472
rect 13145 3366 13179 3400
rect 13275 3438 13309 3472
rect 13275 3366 13309 3400
rect 13405 3438 13439 3472
rect 13405 3366 13439 3400
rect 13535 3438 13569 3472
rect 13535 3366 13569 3400
rect 13665 3438 13699 3472
rect 13665 3366 13699 3400
rect 13795 3438 13829 3472
rect 13795 3366 13829 3400
rect 13925 3438 13959 3472
rect 13925 3366 13959 3400
rect 14055 3438 14089 3472
rect 14055 3366 14089 3400
rect 14185 3438 14219 3472
rect 14185 3366 14219 3400
rect 14315 3438 14349 3472
rect 14315 3366 14349 3400
rect 14445 3438 14479 3472
rect 14445 3366 14479 3400
rect 14575 3438 14609 3472
rect 14575 3366 14609 3400
rect 14705 3438 14739 3472
rect 14705 3366 14739 3400
rect 14835 3438 14869 3472
rect 14835 3366 14869 3400
rect 14965 3438 14999 3472
rect 14965 3366 14999 3400
rect 15095 3438 15129 3472
rect 15095 3366 15129 3400
rect 24607 3438 24641 3472
rect 24607 3366 24641 3400
rect 24737 3438 24771 3472
rect 24737 3366 24771 3400
rect 24867 3438 24901 3472
rect 24867 3366 24901 3400
rect 24997 3438 25031 3472
rect 24997 3366 25031 3400
rect 25127 3438 25161 3472
rect 25127 3366 25161 3400
rect 25257 3438 25291 3472
rect 25257 3366 25291 3400
rect 25387 3438 25421 3472
rect 25387 3366 25421 3400
rect 25517 3438 25551 3472
rect 25517 3366 25551 3400
rect 25647 3438 25681 3472
rect 25647 3366 25681 3400
rect 25777 3438 25811 3472
rect 25777 3366 25811 3400
rect 25907 3438 25941 3472
rect 25907 3366 25941 3400
rect 26037 3438 26071 3472
rect 26037 3366 26071 3400
rect 26167 3438 26201 3472
rect 26167 3366 26201 3400
rect 26297 3438 26331 3472
rect 26297 3366 26331 3400
rect 26427 3438 26461 3472
rect 26427 3366 26461 3400
rect 26557 3438 26591 3472
rect 26557 3366 26591 3400
rect 26687 3438 26721 3472
rect 26687 3366 26721 3400
rect 13145 2826 13179 2860
rect 13145 2754 13179 2788
rect 13275 2826 13309 2860
rect 13275 2754 13309 2788
rect 13405 2826 13439 2860
rect 13405 2754 13439 2788
rect 13535 2826 13569 2860
rect 13535 2754 13569 2788
rect 13665 2826 13699 2860
rect 13665 2754 13699 2788
rect 13795 2826 13829 2860
rect 13795 2754 13829 2788
rect 13925 2826 13959 2860
rect 13925 2754 13959 2788
rect 14055 2826 14089 2860
rect 14055 2754 14089 2788
rect 14185 2826 14219 2860
rect 14185 2754 14219 2788
rect 14315 2826 14349 2860
rect 14315 2754 14349 2788
rect 14445 2826 14479 2860
rect 14445 2754 14479 2788
rect 14575 2826 14609 2860
rect 14575 2754 14609 2788
rect 14705 2826 14739 2860
rect 14705 2754 14739 2788
rect 14835 2826 14869 2860
rect 14835 2754 14869 2788
rect 14965 2826 14999 2860
rect 14965 2754 14999 2788
rect 15095 2826 15129 2860
rect 15095 2754 15129 2788
rect 15225 2826 15259 2860
rect 15225 2754 15259 2788
rect 15355 2826 15389 2860
rect 15355 2754 15389 2788
rect 15485 2826 15519 2860
rect 15485 2754 15519 2788
rect 24737 2826 24771 2860
rect 24737 2754 24771 2788
rect 24867 2826 24901 2860
rect 24867 2754 24901 2788
rect 24997 2826 25031 2860
rect 24997 2754 25031 2788
rect 25127 2826 25161 2860
rect 25127 2754 25161 2788
rect 25257 2826 25291 2860
rect 25257 2754 25291 2788
rect 25387 2826 25421 2860
rect 25387 2754 25421 2788
rect 25517 2826 25551 2860
rect 25517 2754 25551 2788
rect 25647 2826 25681 2860
rect 25647 2754 25681 2788
rect 25777 2826 25811 2860
rect 25777 2754 25811 2788
rect 25907 2826 25941 2860
rect 25907 2754 25941 2788
rect 26037 2826 26071 2860
rect 26037 2754 26071 2788
rect 26167 2826 26201 2860
rect 26167 2754 26201 2788
rect 26297 2826 26331 2860
rect 26297 2754 26331 2788
rect 26427 2826 26461 2860
rect 26427 2754 26461 2788
rect 26557 2826 26591 2860
rect 26557 2754 26591 2788
rect 26687 2826 26721 2860
rect 26687 2754 26721 2788
rect 26817 2826 26851 2860
rect 26817 2754 26851 2788
rect 26947 2826 26981 2860
rect 26947 2754 26981 2788
rect 27077 2826 27111 2860
rect 27077 2754 27111 2788
rect 13145 2478 13179 2512
rect 13145 2406 13179 2440
rect 13275 2478 13309 2512
rect 13275 2406 13309 2440
rect 13405 2478 13439 2512
rect 13405 2406 13439 2440
rect 13535 2478 13569 2512
rect 13535 2406 13569 2440
rect 13665 2478 13699 2512
rect 13665 2406 13699 2440
rect 13795 2478 13829 2512
rect 13795 2406 13829 2440
rect 13925 2478 13959 2512
rect 13925 2406 13959 2440
rect 14055 2478 14089 2512
rect 14055 2406 14089 2440
rect 14185 2478 14219 2512
rect 14185 2406 14219 2440
rect 14315 2478 14349 2512
rect 14315 2406 14349 2440
rect 14445 2478 14479 2512
rect 14445 2406 14479 2440
rect 14575 2478 14609 2512
rect 14575 2406 14609 2440
rect 14705 2478 14739 2512
rect 14705 2406 14739 2440
rect 14835 2478 14869 2512
rect 14835 2406 14869 2440
rect 14965 2478 14999 2512
rect 14965 2406 14999 2440
rect 15095 2478 15129 2512
rect 15095 2406 15129 2440
rect 15225 2478 15259 2512
rect 15225 2406 15259 2440
rect 15355 2478 15389 2512
rect 15355 2406 15389 2440
rect 24737 2478 24771 2512
rect 24737 2406 24771 2440
rect 24867 2478 24901 2512
rect 24867 2406 24901 2440
rect 24997 2478 25031 2512
rect 24997 2406 25031 2440
rect 25127 2478 25161 2512
rect 25127 2406 25161 2440
rect 25257 2478 25291 2512
rect 25257 2406 25291 2440
rect 25387 2478 25421 2512
rect 25387 2406 25421 2440
rect 25517 2478 25551 2512
rect 25517 2406 25551 2440
rect 25647 2478 25681 2512
rect 25647 2406 25681 2440
rect 25777 2478 25811 2512
rect 25777 2406 25811 2440
rect 25907 2478 25941 2512
rect 25907 2406 25941 2440
rect 26037 2478 26071 2512
rect 26037 2406 26071 2440
rect 26167 2478 26201 2512
rect 26167 2406 26201 2440
rect 26297 2478 26331 2512
rect 26297 2406 26331 2440
rect 26427 2478 26461 2512
rect 26427 2406 26461 2440
rect 26557 2478 26591 2512
rect 26557 2406 26591 2440
rect 26687 2478 26721 2512
rect 26687 2406 26721 2440
rect 26817 2478 26851 2512
rect 26817 2406 26851 2440
rect 26947 2478 26981 2512
rect 26947 2406 26981 2440
<< pdiffc >>
rect 13015 5190 13049 5224
rect 13015 5118 13049 5152
rect 13015 5046 13049 5080
rect 13015 4974 13049 5008
rect 13015 4902 13049 4936
rect 13145 5190 13179 5224
rect 13145 5118 13179 5152
rect 13145 5046 13179 5080
rect 13145 4974 13179 5008
rect 13145 4902 13179 4936
rect 13275 5190 13309 5224
rect 13275 5118 13309 5152
rect 13275 5046 13309 5080
rect 13275 4974 13309 5008
rect 13275 4902 13309 4936
rect 13405 5190 13439 5224
rect 13405 5118 13439 5152
rect 13405 5046 13439 5080
rect 13405 4974 13439 5008
rect 13405 4902 13439 4936
rect 13535 5190 13569 5224
rect 13535 5118 13569 5152
rect 13535 5046 13569 5080
rect 13535 4974 13569 5008
rect 13535 4902 13569 4936
rect 13665 5190 13699 5224
rect 13665 5118 13699 5152
rect 13665 5046 13699 5080
rect 13665 4974 13699 5008
rect 13665 4902 13699 4936
rect 13795 5190 13829 5224
rect 13795 5118 13829 5152
rect 13795 5046 13829 5080
rect 13795 4974 13829 5008
rect 13795 4902 13829 4936
rect 13925 5190 13959 5224
rect 13925 5118 13959 5152
rect 13925 5046 13959 5080
rect 13925 4974 13959 5008
rect 13925 4902 13959 4936
rect 14055 5190 14089 5224
rect 14055 5118 14089 5152
rect 14055 5046 14089 5080
rect 14055 4974 14089 5008
rect 14055 4902 14089 4936
rect 14185 5190 14219 5224
rect 14185 5118 14219 5152
rect 14185 5046 14219 5080
rect 14185 4974 14219 5008
rect 14185 4902 14219 4936
rect 14315 5190 14349 5224
rect 14315 5118 14349 5152
rect 14315 5046 14349 5080
rect 14315 4974 14349 5008
rect 14315 4902 14349 4936
rect 14445 5190 14479 5224
rect 14445 5118 14479 5152
rect 14445 5046 14479 5080
rect 14445 4974 14479 5008
rect 14445 4902 14479 4936
rect 14575 5190 14609 5224
rect 14575 5118 14609 5152
rect 14575 5046 14609 5080
rect 14575 4974 14609 5008
rect 14575 4902 14609 4936
rect 14705 5190 14739 5224
rect 14705 5118 14739 5152
rect 14705 5046 14739 5080
rect 14705 4974 14739 5008
rect 14705 4902 14739 4936
rect 14835 5190 14869 5224
rect 14835 5118 14869 5152
rect 14835 5046 14869 5080
rect 14835 4974 14869 5008
rect 14835 4902 14869 4936
rect 14965 5190 14999 5224
rect 14965 5118 14999 5152
rect 14965 5046 14999 5080
rect 14965 4974 14999 5008
rect 14965 4902 14999 4936
rect 15095 5190 15129 5224
rect 15095 5118 15129 5152
rect 15095 5046 15129 5080
rect 15095 4974 15129 5008
rect 15095 4902 15129 4936
rect 24607 5190 24641 5224
rect 24607 5118 24641 5152
rect 24607 5046 24641 5080
rect 24607 4974 24641 5008
rect 24607 4902 24641 4936
rect 24737 5190 24771 5224
rect 24737 5118 24771 5152
rect 24737 5046 24771 5080
rect 24737 4974 24771 5008
rect 24737 4902 24771 4936
rect 24867 5190 24901 5224
rect 24867 5118 24901 5152
rect 24867 5046 24901 5080
rect 24867 4974 24901 5008
rect 24867 4902 24901 4936
rect 24997 5190 25031 5224
rect 24997 5118 25031 5152
rect 24997 5046 25031 5080
rect 24997 4974 25031 5008
rect 24997 4902 25031 4936
rect 25127 5190 25161 5224
rect 25127 5118 25161 5152
rect 25127 5046 25161 5080
rect 25127 4974 25161 5008
rect 25127 4902 25161 4936
rect 25257 5190 25291 5224
rect 25257 5118 25291 5152
rect 25257 5046 25291 5080
rect 25257 4974 25291 5008
rect 25257 4902 25291 4936
rect 25387 5190 25421 5224
rect 25387 5118 25421 5152
rect 25387 5046 25421 5080
rect 25387 4974 25421 5008
rect 25387 4902 25421 4936
rect 25517 5190 25551 5224
rect 25517 5118 25551 5152
rect 25517 5046 25551 5080
rect 25517 4974 25551 5008
rect 25517 4902 25551 4936
rect 25647 5190 25681 5224
rect 25647 5118 25681 5152
rect 25647 5046 25681 5080
rect 25647 4974 25681 5008
rect 25647 4902 25681 4936
rect 25777 5190 25811 5224
rect 25777 5118 25811 5152
rect 25777 5046 25811 5080
rect 25777 4974 25811 5008
rect 25777 4902 25811 4936
rect 25907 5190 25941 5224
rect 25907 5118 25941 5152
rect 25907 5046 25941 5080
rect 25907 4974 25941 5008
rect 25907 4902 25941 4936
rect 26037 5190 26071 5224
rect 26037 5118 26071 5152
rect 26037 5046 26071 5080
rect 26037 4974 26071 5008
rect 26037 4902 26071 4936
rect 26167 5190 26201 5224
rect 26167 5118 26201 5152
rect 26167 5046 26201 5080
rect 26167 4974 26201 5008
rect 26167 4902 26201 4936
rect 26297 5190 26331 5224
rect 26297 5118 26331 5152
rect 26297 5046 26331 5080
rect 26297 4974 26331 5008
rect 26297 4902 26331 4936
rect 26427 5190 26461 5224
rect 26427 5118 26461 5152
rect 26427 5046 26461 5080
rect 26427 4974 26461 5008
rect 26427 4902 26461 4936
rect 26557 5190 26591 5224
rect 26557 5118 26591 5152
rect 26557 5046 26591 5080
rect 26557 4974 26591 5008
rect 26557 4902 26591 4936
rect 26687 5190 26721 5224
rect 26687 5118 26721 5152
rect 26687 5046 26721 5080
rect 26687 4974 26721 5008
rect 26687 4902 26721 4936
rect 13275 4642 13309 4676
rect 13275 4570 13309 4604
rect 13275 4498 13309 4532
rect 13275 4426 13309 4460
rect 13275 4354 13309 4388
rect 13405 4642 13439 4676
rect 13405 4570 13439 4604
rect 13405 4498 13439 4532
rect 13405 4426 13439 4460
rect 13405 4354 13439 4388
rect 13665 4642 13699 4676
rect 13665 4570 13699 4604
rect 13665 4498 13699 4532
rect 13665 4426 13699 4460
rect 13665 4354 13699 4388
rect 13795 4642 13829 4676
rect 13795 4570 13829 4604
rect 13795 4498 13829 4532
rect 13795 4426 13829 4460
rect 13795 4354 13829 4388
rect 14055 4642 14089 4676
rect 14055 4570 14089 4604
rect 14055 4498 14089 4532
rect 14055 4426 14089 4460
rect 14055 4354 14089 4388
rect 14185 4642 14219 4676
rect 14185 4570 14219 4604
rect 14185 4498 14219 4532
rect 14185 4426 14219 4460
rect 14185 4354 14219 4388
rect 14445 4642 14479 4676
rect 14445 4570 14479 4604
rect 14445 4498 14479 4532
rect 14445 4426 14479 4460
rect 14445 4354 14479 4388
rect 14575 4642 14609 4676
rect 14575 4570 14609 4604
rect 14575 4498 14609 4532
rect 14575 4426 14609 4460
rect 14575 4354 14609 4388
rect 14835 4642 14869 4676
rect 14835 4570 14869 4604
rect 14835 4498 14869 4532
rect 14835 4426 14869 4460
rect 14835 4354 14869 4388
rect 14965 4642 14999 4676
rect 14965 4570 14999 4604
rect 14965 4498 14999 4532
rect 14965 4426 14999 4460
rect 14965 4354 14999 4388
rect 15209 4642 15243 4676
rect 15209 4570 15243 4604
rect 15209 4498 15243 4532
rect 15209 4426 15243 4460
rect 15209 4354 15243 4388
rect 15299 4642 15333 4676
rect 15299 4570 15333 4604
rect 15299 4498 15333 4532
rect 15299 4426 15333 4460
rect 15299 4354 15333 4388
rect 15389 4642 15423 4676
rect 15389 4570 15423 4604
rect 15389 4498 15423 4532
rect 15389 4426 15423 4460
rect 15389 4354 15423 4388
rect 15479 4642 15513 4676
rect 15479 4570 15513 4604
rect 15479 4498 15513 4532
rect 15479 4426 15513 4460
rect 15479 4354 15513 4388
rect 15569 4642 15603 4676
rect 15569 4570 15603 4604
rect 15569 4498 15603 4532
rect 15569 4426 15603 4460
rect 15569 4354 15603 4388
rect 24867 4642 24901 4676
rect 24867 4570 24901 4604
rect 24867 4498 24901 4532
rect 24867 4426 24901 4460
rect 24867 4354 24901 4388
rect 24997 4642 25031 4676
rect 24997 4570 25031 4604
rect 24997 4498 25031 4532
rect 24997 4426 25031 4460
rect 24997 4354 25031 4388
rect 25257 4642 25291 4676
rect 25257 4570 25291 4604
rect 25257 4498 25291 4532
rect 25257 4426 25291 4460
rect 25257 4354 25291 4388
rect 25387 4642 25421 4676
rect 25387 4570 25421 4604
rect 25387 4498 25421 4532
rect 25387 4426 25421 4460
rect 25387 4354 25421 4388
rect 25647 4642 25681 4676
rect 25647 4570 25681 4604
rect 25647 4498 25681 4532
rect 25647 4426 25681 4460
rect 25647 4354 25681 4388
rect 25777 4642 25811 4676
rect 25777 4570 25811 4604
rect 25777 4498 25811 4532
rect 25777 4426 25811 4460
rect 25777 4354 25811 4388
rect 26037 4642 26071 4676
rect 26037 4570 26071 4604
rect 26037 4498 26071 4532
rect 26037 4426 26071 4460
rect 26037 4354 26071 4388
rect 26167 4642 26201 4676
rect 26167 4570 26201 4604
rect 26167 4498 26201 4532
rect 26167 4426 26201 4460
rect 26167 4354 26201 4388
rect 26427 4642 26461 4676
rect 26427 4570 26461 4604
rect 26427 4498 26461 4532
rect 26427 4426 26461 4460
rect 26427 4354 26461 4388
rect 26557 4642 26591 4676
rect 26557 4570 26591 4604
rect 26557 4498 26591 4532
rect 26557 4426 26591 4460
rect 26557 4354 26591 4388
rect 26801 4642 26835 4676
rect 26801 4570 26835 4604
rect 26801 4498 26835 4532
rect 26801 4426 26835 4460
rect 26801 4354 26835 4388
rect 26891 4642 26925 4676
rect 26891 4570 26925 4604
rect 26891 4498 26925 4532
rect 26891 4426 26925 4460
rect 26891 4354 26925 4388
rect 26981 4642 27015 4676
rect 26981 4570 27015 4604
rect 26981 4498 27015 4532
rect 26981 4426 27015 4460
rect 26981 4354 27015 4388
rect 27071 4642 27105 4676
rect 27071 4570 27105 4604
rect 27071 4498 27105 4532
rect 27071 4426 27105 4460
rect 27071 4354 27105 4388
rect 27161 4642 27195 4676
rect 27161 4570 27195 4604
rect 27161 4498 27195 4532
rect 27161 4426 27195 4460
rect 27161 4354 27195 4388
rect 13275 1838 13309 1872
rect 13275 1766 13309 1800
rect 13275 1694 13309 1728
rect 13275 1622 13309 1656
rect 13275 1550 13309 1584
rect 13405 1838 13439 1872
rect 13405 1766 13439 1800
rect 13405 1694 13439 1728
rect 13405 1622 13439 1656
rect 13405 1550 13439 1584
rect 13665 1838 13699 1872
rect 13665 1766 13699 1800
rect 13665 1694 13699 1728
rect 13665 1622 13699 1656
rect 13665 1550 13699 1584
rect 13795 1838 13829 1872
rect 13795 1766 13829 1800
rect 13795 1694 13829 1728
rect 13795 1622 13829 1656
rect 13795 1550 13829 1584
rect 14055 1838 14089 1872
rect 14055 1766 14089 1800
rect 14055 1694 14089 1728
rect 14055 1622 14089 1656
rect 14055 1550 14089 1584
rect 14185 1838 14219 1872
rect 14185 1766 14219 1800
rect 14185 1694 14219 1728
rect 14185 1622 14219 1656
rect 14185 1550 14219 1584
rect 14445 1838 14479 1872
rect 14445 1766 14479 1800
rect 14445 1694 14479 1728
rect 14445 1622 14479 1656
rect 14445 1550 14479 1584
rect 14575 1838 14609 1872
rect 14575 1766 14609 1800
rect 14575 1694 14609 1728
rect 14575 1622 14609 1656
rect 14575 1550 14609 1584
rect 14835 1838 14869 1872
rect 14835 1766 14869 1800
rect 14835 1694 14869 1728
rect 14835 1622 14869 1656
rect 14835 1550 14869 1584
rect 14965 1838 14999 1872
rect 14965 1766 14999 1800
rect 14965 1694 14999 1728
rect 14965 1622 14999 1656
rect 14965 1550 14999 1584
rect 15225 1838 15259 1872
rect 15225 1766 15259 1800
rect 15225 1694 15259 1728
rect 15225 1622 15259 1656
rect 15225 1550 15259 1584
rect 15355 1838 15389 1872
rect 15355 1766 15389 1800
rect 15355 1694 15389 1728
rect 15355 1622 15389 1656
rect 15355 1550 15389 1584
rect 24867 1838 24901 1872
rect 24867 1766 24901 1800
rect 24867 1694 24901 1728
rect 24867 1622 24901 1656
rect 24867 1550 24901 1584
rect 24997 1838 25031 1872
rect 24997 1766 25031 1800
rect 24997 1694 25031 1728
rect 24997 1622 25031 1656
rect 24997 1550 25031 1584
rect 25257 1838 25291 1872
rect 25257 1766 25291 1800
rect 25257 1694 25291 1728
rect 25257 1622 25291 1656
rect 25257 1550 25291 1584
rect 25387 1838 25421 1872
rect 25387 1766 25421 1800
rect 25387 1694 25421 1728
rect 25387 1622 25421 1656
rect 25387 1550 25421 1584
rect 25647 1838 25681 1872
rect 25647 1766 25681 1800
rect 25647 1694 25681 1728
rect 25647 1622 25681 1656
rect 25647 1550 25681 1584
rect 25777 1838 25811 1872
rect 25777 1766 25811 1800
rect 25777 1694 25811 1728
rect 25777 1622 25811 1656
rect 25777 1550 25811 1584
rect 26037 1838 26071 1872
rect 26037 1766 26071 1800
rect 26037 1694 26071 1728
rect 26037 1622 26071 1656
rect 26037 1550 26071 1584
rect 26167 1838 26201 1872
rect 26167 1766 26201 1800
rect 26167 1694 26201 1728
rect 26167 1622 26201 1656
rect 26167 1550 26201 1584
rect 26427 1838 26461 1872
rect 26427 1766 26461 1800
rect 26427 1694 26461 1728
rect 26427 1622 26461 1656
rect 26427 1550 26461 1584
rect 26557 1838 26591 1872
rect 26557 1766 26591 1800
rect 26557 1694 26591 1728
rect 26557 1622 26591 1656
rect 26557 1550 26591 1584
rect 26817 1838 26851 1872
rect 26817 1766 26851 1800
rect 26817 1694 26851 1728
rect 26817 1622 26851 1656
rect 26817 1550 26851 1584
rect 26947 1838 26981 1872
rect 26947 1766 26981 1800
rect 26947 1694 26981 1728
rect 26947 1622 26981 1656
rect 26947 1550 26981 1584
rect 13145 1290 13179 1324
rect 13145 1218 13179 1252
rect 13145 1146 13179 1180
rect 13145 1074 13179 1108
rect 13145 1002 13179 1036
rect 13275 1290 13309 1324
rect 13275 1218 13309 1252
rect 13275 1146 13309 1180
rect 13275 1074 13309 1108
rect 13275 1002 13309 1036
rect 13405 1290 13439 1324
rect 13405 1218 13439 1252
rect 13405 1146 13439 1180
rect 13405 1074 13439 1108
rect 13405 1002 13439 1036
rect 13535 1290 13569 1324
rect 13535 1218 13569 1252
rect 13535 1146 13569 1180
rect 13535 1074 13569 1108
rect 13535 1002 13569 1036
rect 13665 1290 13699 1324
rect 13665 1218 13699 1252
rect 13665 1146 13699 1180
rect 13665 1074 13699 1108
rect 13665 1002 13699 1036
rect 13795 1290 13829 1324
rect 13795 1218 13829 1252
rect 13795 1146 13829 1180
rect 13795 1074 13829 1108
rect 13795 1002 13829 1036
rect 13925 1290 13959 1324
rect 13925 1218 13959 1252
rect 13925 1146 13959 1180
rect 13925 1074 13959 1108
rect 13925 1002 13959 1036
rect 14055 1290 14089 1324
rect 14055 1218 14089 1252
rect 14055 1146 14089 1180
rect 14055 1074 14089 1108
rect 14055 1002 14089 1036
rect 14185 1290 14219 1324
rect 14185 1218 14219 1252
rect 14185 1146 14219 1180
rect 14185 1074 14219 1108
rect 14185 1002 14219 1036
rect 14315 1290 14349 1324
rect 14315 1218 14349 1252
rect 14315 1146 14349 1180
rect 14315 1074 14349 1108
rect 14315 1002 14349 1036
rect 14445 1290 14479 1324
rect 14445 1218 14479 1252
rect 14445 1146 14479 1180
rect 14445 1074 14479 1108
rect 14445 1002 14479 1036
rect 14575 1290 14609 1324
rect 14575 1218 14609 1252
rect 14575 1146 14609 1180
rect 14575 1074 14609 1108
rect 14575 1002 14609 1036
rect 14705 1290 14739 1324
rect 14705 1218 14739 1252
rect 14705 1146 14739 1180
rect 14705 1074 14739 1108
rect 14705 1002 14739 1036
rect 14835 1290 14869 1324
rect 14835 1218 14869 1252
rect 14835 1146 14869 1180
rect 14835 1074 14869 1108
rect 14835 1002 14869 1036
rect 14965 1290 14999 1324
rect 14965 1218 14999 1252
rect 14965 1146 14999 1180
rect 14965 1074 14999 1108
rect 14965 1002 14999 1036
rect 15095 1290 15129 1324
rect 15095 1218 15129 1252
rect 15095 1146 15129 1180
rect 15095 1074 15129 1108
rect 15095 1002 15129 1036
rect 15225 1290 15259 1324
rect 15225 1218 15259 1252
rect 15225 1146 15259 1180
rect 15225 1074 15259 1108
rect 15225 1002 15259 1036
rect 15355 1290 15389 1324
rect 15355 1218 15389 1252
rect 15355 1146 15389 1180
rect 15355 1074 15389 1108
rect 15355 1002 15389 1036
rect 15485 1290 15519 1324
rect 15485 1218 15519 1252
rect 15485 1146 15519 1180
rect 15485 1074 15519 1108
rect 15485 1002 15519 1036
rect 24737 1290 24771 1324
rect 24737 1218 24771 1252
rect 24737 1146 24771 1180
rect 24737 1074 24771 1108
rect 24737 1002 24771 1036
rect 24867 1290 24901 1324
rect 24867 1218 24901 1252
rect 24867 1146 24901 1180
rect 24867 1074 24901 1108
rect 24867 1002 24901 1036
rect 24997 1290 25031 1324
rect 24997 1218 25031 1252
rect 24997 1146 25031 1180
rect 24997 1074 25031 1108
rect 24997 1002 25031 1036
rect 25127 1290 25161 1324
rect 25127 1218 25161 1252
rect 25127 1146 25161 1180
rect 25127 1074 25161 1108
rect 25127 1002 25161 1036
rect 25257 1290 25291 1324
rect 25257 1218 25291 1252
rect 25257 1146 25291 1180
rect 25257 1074 25291 1108
rect 25257 1002 25291 1036
rect 25387 1290 25421 1324
rect 25387 1218 25421 1252
rect 25387 1146 25421 1180
rect 25387 1074 25421 1108
rect 25387 1002 25421 1036
rect 25517 1290 25551 1324
rect 25517 1218 25551 1252
rect 25517 1146 25551 1180
rect 25517 1074 25551 1108
rect 25517 1002 25551 1036
rect 25647 1290 25681 1324
rect 25647 1218 25681 1252
rect 25647 1146 25681 1180
rect 25647 1074 25681 1108
rect 25647 1002 25681 1036
rect 25777 1290 25811 1324
rect 25777 1218 25811 1252
rect 25777 1146 25811 1180
rect 25777 1074 25811 1108
rect 25777 1002 25811 1036
rect 25907 1290 25941 1324
rect 25907 1218 25941 1252
rect 25907 1146 25941 1180
rect 25907 1074 25941 1108
rect 25907 1002 25941 1036
rect 26037 1290 26071 1324
rect 26037 1218 26071 1252
rect 26037 1146 26071 1180
rect 26037 1074 26071 1108
rect 26037 1002 26071 1036
rect 26167 1290 26201 1324
rect 26167 1218 26201 1252
rect 26167 1146 26201 1180
rect 26167 1074 26201 1108
rect 26167 1002 26201 1036
rect 26297 1290 26331 1324
rect 26297 1218 26331 1252
rect 26297 1146 26331 1180
rect 26297 1074 26331 1108
rect 26297 1002 26331 1036
rect 26427 1290 26461 1324
rect 26427 1218 26461 1252
rect 26427 1146 26461 1180
rect 26427 1074 26461 1108
rect 26427 1002 26461 1036
rect 26557 1290 26591 1324
rect 26557 1218 26591 1252
rect 26557 1146 26591 1180
rect 26557 1074 26591 1108
rect 26557 1002 26591 1036
rect 26687 1290 26721 1324
rect 26687 1218 26721 1252
rect 26687 1146 26721 1180
rect 26687 1074 26721 1108
rect 26687 1002 26721 1036
rect 26817 1290 26851 1324
rect 26817 1218 26851 1252
rect 26817 1146 26851 1180
rect 26817 1074 26851 1108
rect 26817 1002 26851 1036
rect 26947 1290 26981 1324
rect 26947 1218 26981 1252
rect 26947 1146 26981 1180
rect 26947 1074 26981 1108
rect 26947 1002 26981 1036
rect 27077 1290 27111 1324
rect 27077 1218 27111 1252
rect 27077 1146 27111 1180
rect 27077 1074 27111 1108
rect 27077 1002 27111 1036
<< psubdiff >>
rect 15287 3579 15527 3591
rect 15287 3545 15322 3579
rect 15356 3545 15390 3579
rect 15424 3545 15458 3579
rect 15492 3545 15527 3579
rect 15287 3533 15527 3545
rect 26879 3579 27119 3591
rect 26879 3545 26914 3579
rect 26948 3545 26982 3579
rect 27016 3545 27050 3579
rect 27084 3545 27119 3579
rect 26879 3533 27119 3545
rect 12998 3130 15502 3153
rect 12998 3096 13022 3130
rect 13056 3096 13104 3130
rect 13138 3096 13204 3130
rect 13238 3096 13272 3130
rect 13306 3096 13340 3130
rect 13374 3096 13408 3130
rect 13442 3096 13476 3130
rect 13510 3096 13594 3130
rect 13628 3096 13662 3130
rect 13696 3096 13730 3130
rect 13764 3096 13798 3130
rect 13832 3096 13866 3130
rect 13900 3096 13984 3130
rect 14018 3096 14052 3130
rect 14086 3096 14120 3130
rect 14154 3096 14188 3130
rect 14222 3096 14256 3130
rect 14290 3096 14374 3130
rect 14408 3096 14442 3130
rect 14476 3096 14510 3130
rect 14544 3096 14578 3130
rect 14612 3096 14646 3130
rect 14680 3096 14764 3130
rect 14798 3096 14832 3130
rect 14866 3096 14900 3130
rect 14934 3096 14968 3130
rect 15002 3096 15036 3130
rect 15070 3096 15154 3130
rect 15188 3096 15222 3130
rect 15256 3096 15290 3130
rect 15324 3096 15358 3130
rect 15392 3096 15426 3130
rect 15460 3096 15502 3130
rect 12998 3073 15502 3096
rect 24590 3130 27094 3153
rect 24590 3096 24614 3130
rect 24648 3096 24696 3130
rect 24730 3096 24796 3130
rect 24830 3096 24864 3130
rect 24898 3096 24932 3130
rect 24966 3096 25000 3130
rect 25034 3096 25068 3130
rect 25102 3096 25186 3130
rect 25220 3096 25254 3130
rect 25288 3096 25322 3130
rect 25356 3096 25390 3130
rect 25424 3096 25458 3130
rect 25492 3096 25576 3130
rect 25610 3096 25644 3130
rect 25678 3096 25712 3130
rect 25746 3096 25780 3130
rect 25814 3096 25848 3130
rect 25882 3096 25966 3130
rect 26000 3096 26034 3130
rect 26068 3096 26102 3130
rect 26136 3096 26170 3130
rect 26204 3096 26238 3130
rect 26272 3096 26356 3130
rect 26390 3096 26424 3130
rect 26458 3096 26492 3130
rect 26526 3096 26560 3130
rect 26594 3096 26628 3130
rect 26662 3096 26746 3130
rect 26780 3096 26814 3130
rect 26848 3096 26882 3130
rect 26916 3096 26950 3130
rect 26984 3096 27018 3130
rect 27052 3096 27094 3130
rect 24590 3073 27094 3096
<< nsubdiff >>
rect 12998 5486 15112 5509
rect 12998 5452 13022 5486
rect 13056 5452 13104 5486
rect 13138 5452 13204 5486
rect 13238 5452 13272 5486
rect 13306 5452 13340 5486
rect 13374 5452 13408 5486
rect 13442 5452 13476 5486
rect 13510 5452 13594 5486
rect 13628 5452 13662 5486
rect 13696 5452 13730 5486
rect 13764 5452 13798 5486
rect 13832 5452 13866 5486
rect 13900 5452 13984 5486
rect 14018 5452 14052 5486
rect 14086 5452 14120 5486
rect 14154 5452 14188 5486
rect 14222 5452 14256 5486
rect 14290 5452 14374 5486
rect 14408 5452 14442 5486
rect 14476 5452 14510 5486
rect 14544 5452 14578 5486
rect 14612 5452 14646 5486
rect 14680 5452 14764 5486
rect 14798 5452 14832 5486
rect 14866 5452 14900 5486
rect 14934 5452 14968 5486
rect 15002 5452 15036 5486
rect 15070 5452 15112 5486
rect 12998 5429 15112 5452
rect 24590 5486 26704 5509
rect 24590 5452 24614 5486
rect 24648 5452 24696 5486
rect 24730 5452 24796 5486
rect 24830 5452 24864 5486
rect 24898 5452 24932 5486
rect 24966 5452 25000 5486
rect 25034 5452 25068 5486
rect 25102 5452 25186 5486
rect 25220 5452 25254 5486
rect 25288 5452 25322 5486
rect 25356 5452 25390 5486
rect 25424 5452 25458 5486
rect 25492 5452 25576 5486
rect 25610 5452 25644 5486
rect 25678 5452 25712 5486
rect 25746 5452 25780 5486
rect 25814 5452 25848 5486
rect 25882 5452 25966 5486
rect 26000 5452 26034 5486
rect 26068 5452 26102 5486
rect 26136 5452 26170 5486
rect 26204 5452 26238 5486
rect 26272 5452 26356 5486
rect 26390 5452 26424 5486
rect 26458 5452 26492 5486
rect 26526 5452 26560 5486
rect 26594 5452 26628 5486
rect 26662 5452 26704 5486
rect 24590 5429 26704 5452
rect 15284 4915 15524 4927
rect 15284 4881 15319 4915
rect 15353 4881 15387 4915
rect 15421 4881 15455 4915
rect 15489 4881 15524 4915
rect 15284 4869 15524 4881
rect 26876 4915 27116 4927
rect 26876 4881 26911 4915
rect 26945 4881 26979 4915
rect 27013 4881 27047 4915
rect 27081 4881 27116 4915
rect 26876 4869 27116 4881
rect 13162 774 15502 797
rect 13162 740 13204 774
rect 13238 740 13272 774
rect 13306 740 13340 774
rect 13374 740 13408 774
rect 13442 740 13476 774
rect 13510 740 13594 774
rect 13628 740 13662 774
rect 13696 740 13730 774
rect 13764 740 13798 774
rect 13832 740 13866 774
rect 13900 740 13984 774
rect 14018 740 14052 774
rect 14086 740 14120 774
rect 14154 740 14188 774
rect 14222 740 14256 774
rect 14290 740 14374 774
rect 14408 740 14442 774
rect 14476 740 14510 774
rect 14544 740 14578 774
rect 14612 740 14646 774
rect 14680 740 14764 774
rect 14798 740 14832 774
rect 14866 740 14900 774
rect 14934 740 14968 774
rect 15002 740 15036 774
rect 15070 740 15154 774
rect 15188 740 15222 774
rect 15256 740 15290 774
rect 15324 740 15358 774
rect 15392 740 15426 774
rect 15460 740 15502 774
rect 13162 717 15502 740
rect 24754 774 27094 797
rect 24754 740 24796 774
rect 24830 740 24864 774
rect 24898 740 24932 774
rect 24966 740 25000 774
rect 25034 740 25068 774
rect 25102 740 25186 774
rect 25220 740 25254 774
rect 25288 740 25322 774
rect 25356 740 25390 774
rect 25424 740 25458 774
rect 25492 740 25576 774
rect 25610 740 25644 774
rect 25678 740 25712 774
rect 25746 740 25780 774
rect 25814 740 25848 774
rect 25882 740 25966 774
rect 26000 740 26034 774
rect 26068 740 26102 774
rect 26136 740 26170 774
rect 26204 740 26238 774
rect 26272 740 26356 774
rect 26390 740 26424 774
rect 26458 740 26492 774
rect 26526 740 26560 774
rect 26594 740 26628 774
rect 26662 740 26746 774
rect 26780 740 26814 774
rect 26848 740 26882 774
rect 26916 740 26950 774
rect 26984 740 27018 774
rect 27052 740 27094 774
rect 24754 717 27094 740
<< psubdiffcont >>
rect 15322 3545 15356 3579
rect 15390 3545 15424 3579
rect 15458 3545 15492 3579
rect 26914 3545 26948 3579
rect 26982 3545 27016 3579
rect 27050 3545 27084 3579
rect 13022 3096 13056 3130
rect 13104 3096 13138 3130
rect 13204 3096 13238 3130
rect 13272 3096 13306 3130
rect 13340 3096 13374 3130
rect 13408 3096 13442 3130
rect 13476 3096 13510 3130
rect 13594 3096 13628 3130
rect 13662 3096 13696 3130
rect 13730 3096 13764 3130
rect 13798 3096 13832 3130
rect 13866 3096 13900 3130
rect 13984 3096 14018 3130
rect 14052 3096 14086 3130
rect 14120 3096 14154 3130
rect 14188 3096 14222 3130
rect 14256 3096 14290 3130
rect 14374 3096 14408 3130
rect 14442 3096 14476 3130
rect 14510 3096 14544 3130
rect 14578 3096 14612 3130
rect 14646 3096 14680 3130
rect 14764 3096 14798 3130
rect 14832 3096 14866 3130
rect 14900 3096 14934 3130
rect 14968 3096 15002 3130
rect 15036 3096 15070 3130
rect 15154 3096 15188 3130
rect 15222 3096 15256 3130
rect 15290 3096 15324 3130
rect 15358 3096 15392 3130
rect 15426 3096 15460 3130
rect 24614 3096 24648 3130
rect 24696 3096 24730 3130
rect 24796 3096 24830 3130
rect 24864 3096 24898 3130
rect 24932 3096 24966 3130
rect 25000 3096 25034 3130
rect 25068 3096 25102 3130
rect 25186 3096 25220 3130
rect 25254 3096 25288 3130
rect 25322 3096 25356 3130
rect 25390 3096 25424 3130
rect 25458 3096 25492 3130
rect 25576 3096 25610 3130
rect 25644 3096 25678 3130
rect 25712 3096 25746 3130
rect 25780 3096 25814 3130
rect 25848 3096 25882 3130
rect 25966 3096 26000 3130
rect 26034 3096 26068 3130
rect 26102 3096 26136 3130
rect 26170 3096 26204 3130
rect 26238 3096 26272 3130
rect 26356 3096 26390 3130
rect 26424 3096 26458 3130
rect 26492 3096 26526 3130
rect 26560 3096 26594 3130
rect 26628 3096 26662 3130
rect 26746 3096 26780 3130
rect 26814 3096 26848 3130
rect 26882 3096 26916 3130
rect 26950 3096 26984 3130
rect 27018 3096 27052 3130
<< nsubdiffcont >>
rect 13022 5452 13056 5486
rect 13104 5452 13138 5486
rect 13204 5452 13238 5486
rect 13272 5452 13306 5486
rect 13340 5452 13374 5486
rect 13408 5452 13442 5486
rect 13476 5452 13510 5486
rect 13594 5452 13628 5486
rect 13662 5452 13696 5486
rect 13730 5452 13764 5486
rect 13798 5452 13832 5486
rect 13866 5452 13900 5486
rect 13984 5452 14018 5486
rect 14052 5452 14086 5486
rect 14120 5452 14154 5486
rect 14188 5452 14222 5486
rect 14256 5452 14290 5486
rect 14374 5452 14408 5486
rect 14442 5452 14476 5486
rect 14510 5452 14544 5486
rect 14578 5452 14612 5486
rect 14646 5452 14680 5486
rect 14764 5452 14798 5486
rect 14832 5452 14866 5486
rect 14900 5452 14934 5486
rect 14968 5452 15002 5486
rect 15036 5452 15070 5486
rect 24614 5452 24648 5486
rect 24696 5452 24730 5486
rect 24796 5452 24830 5486
rect 24864 5452 24898 5486
rect 24932 5452 24966 5486
rect 25000 5452 25034 5486
rect 25068 5452 25102 5486
rect 25186 5452 25220 5486
rect 25254 5452 25288 5486
rect 25322 5452 25356 5486
rect 25390 5452 25424 5486
rect 25458 5452 25492 5486
rect 25576 5452 25610 5486
rect 25644 5452 25678 5486
rect 25712 5452 25746 5486
rect 25780 5452 25814 5486
rect 25848 5452 25882 5486
rect 25966 5452 26000 5486
rect 26034 5452 26068 5486
rect 26102 5452 26136 5486
rect 26170 5452 26204 5486
rect 26238 5452 26272 5486
rect 26356 5452 26390 5486
rect 26424 5452 26458 5486
rect 26492 5452 26526 5486
rect 26560 5452 26594 5486
rect 26628 5452 26662 5486
rect 15319 4881 15353 4915
rect 15387 4881 15421 4915
rect 15455 4881 15489 4915
rect 26911 4881 26945 4915
rect 26979 4881 27013 4915
rect 27047 4881 27081 4915
rect 13204 740 13238 774
rect 13272 740 13306 774
rect 13340 740 13374 774
rect 13408 740 13442 774
rect 13476 740 13510 774
rect 13594 740 13628 774
rect 13662 740 13696 774
rect 13730 740 13764 774
rect 13798 740 13832 774
rect 13866 740 13900 774
rect 13984 740 14018 774
rect 14052 740 14086 774
rect 14120 740 14154 774
rect 14188 740 14222 774
rect 14256 740 14290 774
rect 14374 740 14408 774
rect 14442 740 14476 774
rect 14510 740 14544 774
rect 14578 740 14612 774
rect 14646 740 14680 774
rect 14764 740 14798 774
rect 14832 740 14866 774
rect 14900 740 14934 774
rect 14968 740 15002 774
rect 15036 740 15070 774
rect 15154 740 15188 774
rect 15222 740 15256 774
rect 15290 740 15324 774
rect 15358 740 15392 774
rect 15426 740 15460 774
rect 24796 740 24830 774
rect 24864 740 24898 774
rect 24932 740 24966 774
rect 25000 740 25034 774
rect 25068 740 25102 774
rect 25186 740 25220 774
rect 25254 740 25288 774
rect 25322 740 25356 774
rect 25390 740 25424 774
rect 25458 740 25492 774
rect 25576 740 25610 774
rect 25644 740 25678 774
rect 25712 740 25746 774
rect 25780 740 25814 774
rect 25848 740 25882 774
rect 25966 740 26000 774
rect 26034 740 26068 774
rect 26102 740 26136 774
rect 26170 740 26204 774
rect 26238 740 26272 774
rect 26356 740 26390 774
rect 26424 740 26458 774
rect 26492 740 26526 774
rect 26560 740 26594 774
rect 26628 740 26662 774
rect 26746 740 26780 774
rect 26814 740 26848 774
rect 26882 740 26916 774
rect 26950 740 26984 774
rect 27018 740 27052 774
<< poly >>
rect 13062 5353 13132 5369
rect 13062 5319 13080 5353
rect 13114 5319 13132 5353
rect 13062 5263 13132 5319
rect 13192 5353 13262 5369
rect 13192 5319 13210 5353
rect 13244 5319 13262 5353
rect 13192 5263 13262 5319
rect 13322 5353 13392 5369
rect 13322 5319 13340 5353
rect 13374 5319 13392 5353
rect 13322 5263 13392 5319
rect 13452 5353 13522 5369
rect 13452 5319 13470 5353
rect 13504 5319 13522 5353
rect 13452 5263 13522 5319
rect 13582 5353 13652 5369
rect 13582 5319 13600 5353
rect 13634 5319 13652 5353
rect 13582 5263 13652 5319
rect 13712 5353 13782 5369
rect 13712 5319 13730 5353
rect 13764 5319 13782 5353
rect 13712 5263 13782 5319
rect 13842 5353 13912 5369
rect 13842 5319 13860 5353
rect 13894 5319 13912 5353
rect 13842 5263 13912 5319
rect 13972 5353 14042 5369
rect 13972 5319 13990 5353
rect 14024 5319 14042 5353
rect 13972 5263 14042 5319
rect 14102 5353 14172 5369
rect 14102 5319 14120 5353
rect 14154 5319 14172 5353
rect 14102 5263 14172 5319
rect 14232 5353 14302 5369
rect 14232 5319 14250 5353
rect 14284 5319 14302 5353
rect 14232 5263 14302 5319
rect 14362 5353 14432 5369
rect 14362 5319 14380 5353
rect 14414 5319 14432 5353
rect 14362 5263 14432 5319
rect 14492 5353 14562 5369
rect 14492 5319 14510 5353
rect 14544 5319 14562 5353
rect 14492 5263 14562 5319
rect 14622 5353 14692 5369
rect 14622 5319 14640 5353
rect 14674 5319 14692 5353
rect 14622 5263 14692 5319
rect 14752 5353 14822 5369
rect 14752 5319 14770 5353
rect 14804 5319 14822 5353
rect 14752 5263 14822 5319
rect 14882 5353 14952 5369
rect 14882 5319 14900 5353
rect 14934 5319 14952 5353
rect 14882 5263 14952 5319
rect 15012 5353 15082 5369
rect 15012 5319 15030 5353
rect 15064 5319 15082 5353
rect 15012 5263 15082 5319
rect 24654 5353 24724 5369
rect 24654 5319 24672 5353
rect 24706 5319 24724 5353
rect 24654 5263 24724 5319
rect 24784 5353 24854 5369
rect 24784 5319 24802 5353
rect 24836 5319 24854 5353
rect 24784 5263 24854 5319
rect 24914 5353 24984 5369
rect 24914 5319 24932 5353
rect 24966 5319 24984 5353
rect 24914 5263 24984 5319
rect 25044 5353 25114 5369
rect 25044 5319 25062 5353
rect 25096 5319 25114 5353
rect 25044 5263 25114 5319
rect 25174 5353 25244 5369
rect 25174 5319 25192 5353
rect 25226 5319 25244 5353
rect 25174 5263 25244 5319
rect 25304 5353 25374 5369
rect 25304 5319 25322 5353
rect 25356 5319 25374 5353
rect 25304 5263 25374 5319
rect 25434 5353 25504 5369
rect 25434 5319 25452 5353
rect 25486 5319 25504 5353
rect 25434 5263 25504 5319
rect 25564 5353 25634 5369
rect 25564 5319 25582 5353
rect 25616 5319 25634 5353
rect 25564 5263 25634 5319
rect 25694 5353 25764 5369
rect 25694 5319 25712 5353
rect 25746 5319 25764 5353
rect 25694 5263 25764 5319
rect 25824 5353 25894 5369
rect 25824 5319 25842 5353
rect 25876 5319 25894 5353
rect 25824 5263 25894 5319
rect 25954 5353 26024 5369
rect 25954 5319 25972 5353
rect 26006 5319 26024 5353
rect 25954 5263 26024 5319
rect 26084 5353 26154 5369
rect 26084 5319 26102 5353
rect 26136 5319 26154 5353
rect 26084 5263 26154 5319
rect 26214 5353 26284 5369
rect 26214 5319 26232 5353
rect 26266 5319 26284 5353
rect 26214 5263 26284 5319
rect 26344 5353 26414 5369
rect 26344 5319 26362 5353
rect 26396 5319 26414 5353
rect 26344 5263 26414 5319
rect 26474 5353 26544 5369
rect 26474 5319 26492 5353
rect 26526 5319 26544 5353
rect 26474 5263 26544 5319
rect 26604 5353 26674 5369
rect 26604 5319 26622 5353
rect 26656 5319 26674 5353
rect 26604 5263 26674 5319
rect 13062 4823 13132 4863
rect 13192 4823 13262 4863
rect 13322 4823 13392 4863
rect 13452 4823 13522 4863
rect 13582 4823 13652 4863
rect 13712 4823 13782 4863
rect 13842 4823 13912 4863
rect 13972 4823 14042 4863
rect 14102 4823 14172 4863
rect 14232 4823 14302 4863
rect 14362 4823 14432 4863
rect 14492 4823 14562 4863
rect 14622 4823 14692 4863
rect 14752 4823 14822 4863
rect 14882 4823 14952 4863
rect 15012 4823 15082 4863
rect 15346 4824 15556 4834
rect 15346 4790 15404 4824
rect 15438 4790 15472 4824
rect 15506 4790 15556 4824
rect 24654 4823 24724 4863
rect 24784 4823 24854 4863
rect 24914 4823 24984 4863
rect 25044 4823 25114 4863
rect 25174 4823 25244 4863
rect 25304 4823 25374 4863
rect 25434 4823 25504 4863
rect 25564 4823 25634 4863
rect 25694 4823 25764 4863
rect 25824 4823 25894 4863
rect 25954 4823 26024 4863
rect 26084 4823 26154 4863
rect 26214 4823 26284 4863
rect 26344 4823 26414 4863
rect 26474 4823 26544 4863
rect 26604 4823 26674 4863
rect 26938 4824 27148 4834
rect 15346 4780 15556 4790
rect 13322 4715 13392 4755
rect 13712 4715 13782 4755
rect 14102 4715 14172 4755
rect 14492 4715 14562 4755
rect 14882 4715 14952 4755
rect 15256 4715 15286 4755
rect 15346 4715 15376 4780
rect 15436 4715 15466 4780
rect 15526 4715 15556 4780
rect 26938 4790 26996 4824
rect 27030 4790 27064 4824
rect 27098 4790 27148 4824
rect 26938 4780 27148 4790
rect 24914 4715 24984 4755
rect 25304 4715 25374 4755
rect 25694 4715 25764 4755
rect 26084 4715 26154 4755
rect 26474 4715 26544 4755
rect 26848 4715 26878 4755
rect 26938 4715 26968 4780
rect 27028 4715 27058 4780
rect 27118 4715 27148 4780
rect 13322 4123 13392 4315
rect 13712 4123 13782 4315
rect 14102 4123 14172 4315
rect 14492 4123 14562 4315
rect 14882 4123 14952 4315
rect 13228 4108 13392 4123
rect 13228 4074 13244 4108
rect 13278 4074 13392 4108
rect 13228 4059 13392 4074
rect 13618 4108 13782 4123
rect 13618 4074 13634 4108
rect 13668 4074 13782 4108
rect 13618 4059 13782 4074
rect 14008 4108 14172 4123
rect 14008 4074 14024 4108
rect 14058 4074 14172 4108
rect 14008 4059 14172 4074
rect 14398 4108 14562 4123
rect 14398 4074 14414 4108
rect 14448 4074 14562 4108
rect 14398 4059 14562 4074
rect 14788 4108 14952 4123
rect 15256 4118 15286 4315
rect 14788 4074 14804 4108
rect 14838 4074 14952 4108
rect 14788 4059 14952 4074
rect 15233 4108 15299 4118
rect 15233 4074 15249 4108
rect 15283 4074 15299 4108
rect 15233 4064 15299 4074
rect 13322 3867 13392 4059
rect 13452 3867 13522 3907
rect 13712 3867 13782 4059
rect 13842 3951 13912 3961
rect 13842 3917 13860 3951
rect 13894 3917 13912 3951
rect 13842 3867 13912 3917
rect 14102 3867 14172 4059
rect 14232 3867 14302 3907
rect 14492 3867 14562 4059
rect 14622 3951 14692 3961
rect 14622 3917 14640 3951
rect 14674 3917 14692 3951
rect 14622 3867 14692 3917
rect 14882 3867 14952 4059
rect 15012 3867 15082 3907
rect 15256 3867 15286 4064
rect 15346 3867 15376 4315
rect 15436 3867 15466 4315
rect 15526 3867 15556 4315
rect 24914 4123 24984 4315
rect 25304 4123 25374 4315
rect 25694 4123 25764 4315
rect 26084 4123 26154 4315
rect 26474 4123 26544 4315
rect 24820 4108 24984 4123
rect 24820 4074 24836 4108
rect 24870 4074 24984 4108
rect 24820 4059 24984 4074
rect 25210 4108 25374 4123
rect 25210 4074 25226 4108
rect 25260 4074 25374 4108
rect 25210 4059 25374 4074
rect 25600 4108 25764 4123
rect 25600 4074 25616 4108
rect 25650 4074 25764 4108
rect 25600 4059 25764 4074
rect 25990 4108 26154 4123
rect 25990 4074 26006 4108
rect 26040 4074 26154 4108
rect 25990 4059 26154 4074
rect 26380 4108 26544 4123
rect 26848 4118 26878 4315
rect 26380 4074 26396 4108
rect 26430 4074 26544 4108
rect 26380 4059 26544 4074
rect 26825 4108 26891 4118
rect 26825 4074 26841 4108
rect 26875 4074 26891 4108
rect 26825 4064 26891 4074
rect 24914 3867 24984 4059
rect 25044 3867 25114 3907
rect 25304 3867 25374 4059
rect 25434 3951 25504 3961
rect 25434 3917 25452 3951
rect 25486 3917 25504 3951
rect 25434 3867 25504 3917
rect 25694 3867 25764 4059
rect 25824 3867 25894 3907
rect 26084 3867 26154 4059
rect 26214 3951 26284 3961
rect 26214 3917 26232 3951
rect 26266 3917 26284 3951
rect 26214 3867 26284 3917
rect 26474 3867 26544 4059
rect 26604 3867 26674 3907
rect 26848 3867 26878 4064
rect 26938 3867 26968 4315
rect 27028 3867 27058 4315
rect 27118 3867 27148 4315
rect 13322 3627 13392 3667
rect 13062 3519 13132 3559
rect 13192 3519 13262 3559
rect 13322 3519 13392 3559
rect 13452 3519 13522 3667
rect 13712 3627 13782 3667
rect 13842 3627 13912 3667
rect 14102 3627 14172 3667
rect 13582 3519 13652 3559
rect 13712 3519 13782 3559
rect 13842 3519 13912 3559
rect 13972 3519 14042 3559
rect 14102 3519 14172 3559
rect 14232 3519 14302 3667
rect 14492 3627 14562 3667
rect 14622 3627 14692 3667
rect 14882 3627 14952 3667
rect 14362 3519 14432 3559
rect 14492 3519 14562 3559
rect 14622 3519 14692 3559
rect 14752 3519 14822 3559
rect 14882 3519 14952 3559
rect 15012 3519 15082 3667
rect 15256 3627 15286 3667
rect 15346 3627 15376 3667
rect 15436 3627 15466 3667
rect 15526 3627 15556 3667
rect 24914 3627 24984 3667
rect 24654 3519 24724 3559
rect 24784 3519 24854 3559
rect 24914 3519 24984 3559
rect 25044 3519 25114 3667
rect 25304 3627 25374 3667
rect 25434 3627 25504 3667
rect 25694 3627 25764 3667
rect 25174 3519 25244 3559
rect 25304 3519 25374 3559
rect 25434 3519 25504 3559
rect 25564 3519 25634 3559
rect 25694 3519 25764 3559
rect 25824 3519 25894 3667
rect 26084 3627 26154 3667
rect 26214 3627 26284 3667
rect 26474 3627 26544 3667
rect 25954 3519 26024 3559
rect 26084 3519 26154 3559
rect 26214 3519 26284 3559
rect 26344 3519 26414 3559
rect 26474 3519 26544 3559
rect 26604 3519 26674 3667
rect 26848 3627 26878 3667
rect 26938 3627 26968 3667
rect 27028 3627 27058 3667
rect 27118 3627 27148 3667
rect 13062 3279 13132 3319
rect 12996 3263 13132 3279
rect 12996 3229 13012 3263
rect 13046 3229 13132 3263
rect 12996 3213 13132 3229
rect 13192 3263 13262 3319
rect 13192 3229 13210 3263
rect 13244 3229 13262 3263
rect 13192 3213 13262 3229
rect 13322 3263 13392 3319
rect 13322 3229 13340 3263
rect 13374 3229 13392 3263
rect 13322 3213 13392 3229
rect 13452 3263 13522 3319
rect 13452 3229 13470 3263
rect 13504 3229 13522 3263
rect 13452 3213 13522 3229
rect 13582 3263 13652 3319
rect 13582 3229 13600 3263
rect 13634 3229 13652 3263
rect 13582 3213 13652 3229
rect 13712 3263 13782 3319
rect 13712 3229 13730 3263
rect 13764 3229 13782 3263
rect 13712 3213 13782 3229
rect 13842 3263 13912 3319
rect 13842 3229 13860 3263
rect 13894 3229 13912 3263
rect 13842 3213 13912 3229
rect 13972 3263 14042 3319
rect 13972 3229 13990 3263
rect 14024 3229 14042 3263
rect 13972 3213 14042 3229
rect 14102 3263 14172 3319
rect 14102 3229 14120 3263
rect 14154 3229 14172 3263
rect 14102 3213 14172 3229
rect 14232 3263 14302 3319
rect 14232 3229 14250 3263
rect 14284 3229 14302 3263
rect 14232 3213 14302 3229
rect 14362 3263 14432 3319
rect 14362 3229 14380 3263
rect 14414 3229 14432 3263
rect 14362 3213 14432 3229
rect 14492 3263 14562 3319
rect 14492 3229 14510 3263
rect 14544 3229 14562 3263
rect 14492 3213 14562 3229
rect 14622 3263 14692 3319
rect 14622 3229 14640 3263
rect 14674 3229 14692 3263
rect 14622 3213 14692 3229
rect 14752 3263 14822 3319
rect 14752 3229 14770 3263
rect 14804 3229 14822 3263
rect 14752 3213 14822 3229
rect 14882 3263 14952 3319
rect 14882 3229 14900 3263
rect 14934 3229 14952 3263
rect 14882 3213 14952 3229
rect 15012 3263 15082 3319
rect 24654 3279 24724 3319
rect 15012 3229 15030 3263
rect 15064 3229 15082 3263
rect 15012 3213 15082 3229
rect 24588 3263 24724 3279
rect 24588 3229 24604 3263
rect 24638 3229 24724 3263
rect 24588 3213 24724 3229
rect 24784 3263 24854 3319
rect 24784 3229 24802 3263
rect 24836 3229 24854 3263
rect 24784 3213 24854 3229
rect 24914 3263 24984 3319
rect 24914 3229 24932 3263
rect 24966 3229 24984 3263
rect 24914 3213 24984 3229
rect 25044 3263 25114 3319
rect 25044 3229 25062 3263
rect 25096 3229 25114 3263
rect 25044 3213 25114 3229
rect 25174 3263 25244 3319
rect 25174 3229 25192 3263
rect 25226 3229 25244 3263
rect 25174 3213 25244 3229
rect 25304 3263 25374 3319
rect 25304 3229 25322 3263
rect 25356 3229 25374 3263
rect 25304 3213 25374 3229
rect 25434 3263 25504 3319
rect 25434 3229 25452 3263
rect 25486 3229 25504 3263
rect 25434 3213 25504 3229
rect 25564 3263 25634 3319
rect 25564 3229 25582 3263
rect 25616 3229 25634 3263
rect 25564 3213 25634 3229
rect 25694 3263 25764 3319
rect 25694 3229 25712 3263
rect 25746 3229 25764 3263
rect 25694 3213 25764 3229
rect 25824 3263 25894 3319
rect 25824 3229 25842 3263
rect 25876 3229 25894 3263
rect 25824 3213 25894 3229
rect 25954 3263 26024 3319
rect 25954 3229 25972 3263
rect 26006 3229 26024 3263
rect 25954 3213 26024 3229
rect 26084 3263 26154 3319
rect 26084 3229 26102 3263
rect 26136 3229 26154 3263
rect 26084 3213 26154 3229
rect 26214 3263 26284 3319
rect 26214 3229 26232 3263
rect 26266 3229 26284 3263
rect 26214 3213 26284 3229
rect 26344 3263 26414 3319
rect 26344 3229 26362 3263
rect 26396 3229 26414 3263
rect 26344 3213 26414 3229
rect 26474 3263 26544 3319
rect 26474 3229 26492 3263
rect 26526 3229 26544 3263
rect 26474 3213 26544 3229
rect 26604 3263 26674 3319
rect 26604 3229 26622 3263
rect 26656 3229 26674 3263
rect 26604 3213 26674 3229
rect 13192 2997 13262 3013
rect 13192 2963 13210 2997
rect 13244 2963 13262 2997
rect 13192 2907 13262 2963
rect 13322 2997 13392 3013
rect 13322 2963 13340 2997
rect 13374 2963 13392 2997
rect 13322 2907 13392 2963
rect 13452 2997 13522 3013
rect 13452 2963 13470 2997
rect 13504 2963 13522 2997
rect 13452 2907 13522 2963
rect 13582 2997 13652 3013
rect 13582 2963 13600 2997
rect 13634 2963 13652 2997
rect 13582 2907 13652 2963
rect 13712 2997 13782 3013
rect 13712 2963 13730 2997
rect 13764 2963 13782 2997
rect 13712 2907 13782 2963
rect 13842 2997 13912 3013
rect 13842 2963 13860 2997
rect 13894 2963 13912 2997
rect 13842 2907 13912 2963
rect 13972 2997 14042 3013
rect 13972 2963 13990 2997
rect 14024 2963 14042 2997
rect 13972 2907 14042 2963
rect 14102 2997 14172 3013
rect 14102 2963 14120 2997
rect 14154 2963 14172 2997
rect 14102 2907 14172 2963
rect 14232 2997 14302 3013
rect 14232 2963 14250 2997
rect 14284 2963 14302 2997
rect 14232 2907 14302 2963
rect 14362 2997 14432 3013
rect 14362 2963 14380 2997
rect 14414 2963 14432 2997
rect 14362 2907 14432 2963
rect 14492 2997 14562 3013
rect 14492 2963 14510 2997
rect 14544 2963 14562 2997
rect 14492 2907 14562 2963
rect 14622 2997 14692 3013
rect 14622 2963 14640 2997
rect 14674 2963 14692 2997
rect 14622 2907 14692 2963
rect 14752 2997 14822 3013
rect 14752 2963 14770 2997
rect 14804 2963 14822 2997
rect 14752 2907 14822 2963
rect 14882 2997 14952 3013
rect 14882 2963 14900 2997
rect 14934 2963 14952 2997
rect 14882 2907 14952 2963
rect 15012 2997 15082 3013
rect 15012 2963 15030 2997
rect 15064 2963 15082 2997
rect 15012 2907 15082 2963
rect 15142 2997 15212 3013
rect 15142 2963 15160 2997
rect 15194 2963 15212 2997
rect 15142 2907 15212 2963
rect 15272 2997 15342 3013
rect 15272 2963 15290 2997
rect 15324 2963 15342 2997
rect 15272 2907 15342 2963
rect 15402 2997 15472 3013
rect 15402 2963 15420 2997
rect 15454 2963 15472 2997
rect 15402 2907 15472 2963
rect 24784 2997 24854 3013
rect 24784 2963 24802 2997
rect 24836 2963 24854 2997
rect 24784 2907 24854 2963
rect 24914 2997 24984 3013
rect 24914 2963 24932 2997
rect 24966 2963 24984 2997
rect 24914 2907 24984 2963
rect 25044 2997 25114 3013
rect 25044 2963 25062 2997
rect 25096 2963 25114 2997
rect 25044 2907 25114 2963
rect 25174 2997 25244 3013
rect 25174 2963 25192 2997
rect 25226 2963 25244 2997
rect 25174 2907 25244 2963
rect 25304 2997 25374 3013
rect 25304 2963 25322 2997
rect 25356 2963 25374 2997
rect 25304 2907 25374 2963
rect 25434 2997 25504 3013
rect 25434 2963 25452 2997
rect 25486 2963 25504 2997
rect 25434 2907 25504 2963
rect 25564 2997 25634 3013
rect 25564 2963 25582 2997
rect 25616 2963 25634 2997
rect 25564 2907 25634 2963
rect 25694 2997 25764 3013
rect 25694 2963 25712 2997
rect 25746 2963 25764 2997
rect 25694 2907 25764 2963
rect 25824 2997 25894 3013
rect 25824 2963 25842 2997
rect 25876 2963 25894 2997
rect 25824 2907 25894 2963
rect 25954 2997 26024 3013
rect 25954 2963 25972 2997
rect 26006 2963 26024 2997
rect 25954 2907 26024 2963
rect 26084 2997 26154 3013
rect 26084 2963 26102 2997
rect 26136 2963 26154 2997
rect 26084 2907 26154 2963
rect 26214 2997 26284 3013
rect 26214 2963 26232 2997
rect 26266 2963 26284 2997
rect 26214 2907 26284 2963
rect 26344 2997 26414 3013
rect 26344 2963 26362 2997
rect 26396 2963 26414 2997
rect 26344 2907 26414 2963
rect 26474 2997 26544 3013
rect 26474 2963 26492 2997
rect 26526 2963 26544 2997
rect 26474 2907 26544 2963
rect 26604 2997 26674 3013
rect 26604 2963 26622 2997
rect 26656 2963 26674 2997
rect 26604 2907 26674 2963
rect 26734 2997 26804 3013
rect 26734 2963 26752 2997
rect 26786 2963 26804 2997
rect 26734 2907 26804 2963
rect 26864 2997 26934 3013
rect 26864 2963 26882 2997
rect 26916 2963 26934 2997
rect 26864 2907 26934 2963
rect 26994 2997 27064 3013
rect 26994 2963 27012 2997
rect 27046 2963 27064 2997
rect 26994 2907 27064 2963
rect 13192 2667 13262 2707
rect 13322 2667 13392 2707
rect 13452 2667 13522 2707
rect 13582 2667 13652 2707
rect 13712 2667 13782 2707
rect 13842 2667 13912 2707
rect 13192 2559 13262 2599
rect 13322 2559 13392 2599
rect 13582 2559 13652 2599
rect 13712 2559 13782 2599
rect 13972 2559 14042 2707
rect 14102 2667 14172 2707
rect 14232 2667 14302 2707
rect 14362 2667 14432 2707
rect 14492 2667 14562 2707
rect 14622 2667 14692 2707
rect 14102 2559 14172 2599
rect 14362 2559 14432 2599
rect 14492 2559 14562 2599
rect 14752 2559 14822 2707
rect 14882 2667 14952 2707
rect 15012 2667 15082 2707
rect 15142 2667 15212 2707
rect 15272 2667 15342 2707
rect 15402 2667 15472 2707
rect 24784 2667 24854 2707
rect 24914 2667 24984 2707
rect 25044 2667 25114 2707
rect 25174 2667 25244 2707
rect 25304 2667 25374 2707
rect 25434 2667 25504 2707
rect 14882 2559 14952 2599
rect 15142 2559 15212 2599
rect 15272 2559 15342 2599
rect 24784 2559 24854 2599
rect 24914 2559 24984 2599
rect 25174 2559 25244 2599
rect 25304 2559 25374 2599
rect 25564 2559 25634 2707
rect 25694 2667 25764 2707
rect 25824 2667 25894 2707
rect 25954 2667 26024 2707
rect 26084 2667 26154 2707
rect 26214 2667 26284 2707
rect 25694 2559 25764 2599
rect 25954 2559 26024 2599
rect 26084 2559 26154 2599
rect 26344 2559 26414 2707
rect 26474 2667 26544 2707
rect 26604 2667 26674 2707
rect 26734 2667 26804 2707
rect 26864 2667 26934 2707
rect 26994 2667 27064 2707
rect 26474 2559 26544 2599
rect 26734 2559 26804 2599
rect 26864 2559 26934 2599
rect 13192 2309 13262 2359
rect 13192 2275 13210 2309
rect 13244 2275 13262 2309
rect 13192 2265 13262 2275
rect 13322 2167 13392 2359
rect 13582 2309 13652 2359
rect 13582 2275 13600 2309
rect 13634 2275 13652 2309
rect 13582 2265 13652 2275
rect 13712 2167 13782 2359
rect 13972 2319 14042 2359
rect 14102 2167 14172 2359
rect 14362 2309 14432 2359
rect 14362 2275 14380 2309
rect 14414 2275 14432 2309
rect 14362 2265 14432 2275
rect 14492 2167 14562 2359
rect 14752 2319 14822 2359
rect 14882 2167 14952 2359
rect 15142 2309 15212 2359
rect 15142 2275 15160 2309
rect 15194 2275 15212 2309
rect 15142 2265 15212 2275
rect 15272 2167 15342 2359
rect 24784 2309 24854 2359
rect 24784 2275 24802 2309
rect 24836 2275 24854 2309
rect 24784 2265 24854 2275
rect 24914 2167 24984 2359
rect 25174 2309 25244 2359
rect 25174 2275 25192 2309
rect 25226 2275 25244 2309
rect 25174 2265 25244 2275
rect 25304 2167 25374 2359
rect 25564 2319 25634 2359
rect 25694 2167 25764 2359
rect 25954 2309 26024 2359
rect 25954 2275 25972 2309
rect 26006 2275 26024 2309
rect 25954 2265 26024 2275
rect 26084 2167 26154 2359
rect 26344 2319 26414 2359
rect 26474 2167 26544 2359
rect 26734 2309 26804 2359
rect 26734 2275 26752 2309
rect 26786 2275 26804 2309
rect 26734 2265 26804 2275
rect 26864 2167 26934 2359
rect 13322 2152 13486 2167
rect 13322 2118 13436 2152
rect 13470 2118 13486 2152
rect 13322 2103 13486 2118
rect 13712 2152 13876 2167
rect 13712 2118 13826 2152
rect 13860 2118 13876 2152
rect 13712 2103 13876 2118
rect 14102 2152 14266 2167
rect 14102 2118 14216 2152
rect 14250 2118 14266 2152
rect 14102 2103 14266 2118
rect 14492 2152 14656 2167
rect 14492 2118 14606 2152
rect 14640 2118 14656 2152
rect 14492 2103 14656 2118
rect 14882 2152 15046 2167
rect 14882 2118 14996 2152
rect 15030 2118 15046 2152
rect 14882 2103 15046 2118
rect 15272 2152 15436 2167
rect 15272 2118 15386 2152
rect 15420 2118 15436 2152
rect 15272 2103 15436 2118
rect 24914 2152 25078 2167
rect 24914 2118 25028 2152
rect 25062 2118 25078 2152
rect 24914 2103 25078 2118
rect 25304 2152 25468 2167
rect 25304 2118 25418 2152
rect 25452 2118 25468 2152
rect 25304 2103 25468 2118
rect 25694 2152 25858 2167
rect 25694 2118 25808 2152
rect 25842 2118 25858 2152
rect 25694 2103 25858 2118
rect 26084 2152 26248 2167
rect 26084 2118 26198 2152
rect 26232 2118 26248 2152
rect 26084 2103 26248 2118
rect 26474 2152 26638 2167
rect 26474 2118 26588 2152
rect 26622 2118 26638 2152
rect 26474 2103 26638 2118
rect 26864 2152 27028 2167
rect 26864 2118 26978 2152
rect 27012 2118 27028 2152
rect 26864 2103 27028 2118
rect 13322 1911 13392 2103
rect 13712 1911 13782 2103
rect 14102 1911 14172 2103
rect 14492 1911 14562 2103
rect 14882 1911 14952 2103
rect 15272 1911 15342 2103
rect 24914 1911 24984 2103
rect 25304 1911 25374 2103
rect 25694 1911 25764 2103
rect 26084 1911 26154 2103
rect 26474 1911 26544 2103
rect 26864 1911 26934 2103
rect 13322 1471 13392 1511
rect 13712 1471 13782 1511
rect 14102 1471 14172 1511
rect 14492 1471 14562 1511
rect 14882 1471 14952 1511
rect 15272 1471 15342 1511
rect 24914 1471 24984 1511
rect 25304 1471 25374 1511
rect 25694 1471 25764 1511
rect 26084 1471 26154 1511
rect 26474 1471 26544 1511
rect 26864 1471 26934 1511
rect 13192 1363 13262 1403
rect 13322 1363 13392 1403
rect 13452 1363 13522 1403
rect 13582 1363 13652 1403
rect 13712 1363 13782 1403
rect 13842 1363 13912 1403
rect 13972 1363 14042 1403
rect 14102 1363 14172 1403
rect 14232 1363 14302 1403
rect 14362 1363 14432 1403
rect 14492 1363 14562 1403
rect 14622 1363 14692 1403
rect 14752 1363 14822 1403
rect 14882 1363 14952 1403
rect 15012 1363 15082 1403
rect 15142 1363 15212 1403
rect 15272 1363 15342 1403
rect 15402 1363 15472 1403
rect 24784 1363 24854 1403
rect 24914 1363 24984 1403
rect 25044 1363 25114 1403
rect 25174 1363 25244 1403
rect 25304 1363 25374 1403
rect 25434 1363 25504 1403
rect 25564 1363 25634 1403
rect 25694 1363 25764 1403
rect 25824 1363 25894 1403
rect 25954 1363 26024 1403
rect 26084 1363 26154 1403
rect 26214 1363 26284 1403
rect 26344 1363 26414 1403
rect 26474 1363 26544 1403
rect 26604 1363 26674 1403
rect 26734 1363 26804 1403
rect 26864 1363 26934 1403
rect 26994 1363 27064 1403
rect 13192 907 13262 963
rect 13192 873 13210 907
rect 13244 873 13262 907
rect 13192 857 13262 873
rect 13322 907 13392 963
rect 13322 873 13340 907
rect 13374 873 13392 907
rect 13322 857 13392 873
rect 13452 907 13522 963
rect 13452 873 13470 907
rect 13504 873 13522 907
rect 13452 857 13522 873
rect 13582 907 13652 963
rect 13582 873 13600 907
rect 13634 873 13652 907
rect 13582 857 13652 873
rect 13712 907 13782 963
rect 13712 873 13730 907
rect 13764 873 13782 907
rect 13712 857 13782 873
rect 13842 907 13912 963
rect 13842 873 13860 907
rect 13894 873 13912 907
rect 13842 857 13912 873
rect 13972 907 14042 963
rect 13972 873 13990 907
rect 14024 873 14042 907
rect 13972 857 14042 873
rect 14102 907 14172 963
rect 14102 873 14120 907
rect 14154 873 14172 907
rect 14102 857 14172 873
rect 14232 907 14302 963
rect 14232 873 14250 907
rect 14284 873 14302 907
rect 14232 857 14302 873
rect 14362 907 14432 963
rect 14362 873 14380 907
rect 14414 873 14432 907
rect 14362 857 14432 873
rect 14492 907 14562 963
rect 14492 873 14510 907
rect 14544 873 14562 907
rect 14492 857 14562 873
rect 14622 907 14692 963
rect 14622 873 14640 907
rect 14674 873 14692 907
rect 14622 857 14692 873
rect 14752 907 14822 963
rect 14752 873 14770 907
rect 14804 873 14822 907
rect 14752 857 14822 873
rect 14882 907 14952 963
rect 14882 873 14900 907
rect 14934 873 14952 907
rect 14882 857 14952 873
rect 15012 907 15082 963
rect 15012 873 15030 907
rect 15064 873 15082 907
rect 15012 857 15082 873
rect 15142 907 15212 963
rect 15142 873 15160 907
rect 15194 873 15212 907
rect 15142 857 15212 873
rect 15272 907 15342 963
rect 15272 873 15290 907
rect 15324 873 15342 907
rect 15272 857 15342 873
rect 15402 907 15472 963
rect 15402 873 15420 907
rect 15454 873 15472 907
rect 15402 857 15472 873
rect 24784 907 24854 963
rect 24784 873 24802 907
rect 24836 873 24854 907
rect 24784 857 24854 873
rect 24914 907 24984 963
rect 24914 873 24932 907
rect 24966 873 24984 907
rect 24914 857 24984 873
rect 25044 907 25114 963
rect 25044 873 25062 907
rect 25096 873 25114 907
rect 25044 857 25114 873
rect 25174 907 25244 963
rect 25174 873 25192 907
rect 25226 873 25244 907
rect 25174 857 25244 873
rect 25304 907 25374 963
rect 25304 873 25322 907
rect 25356 873 25374 907
rect 25304 857 25374 873
rect 25434 907 25504 963
rect 25434 873 25452 907
rect 25486 873 25504 907
rect 25434 857 25504 873
rect 25564 907 25634 963
rect 25564 873 25582 907
rect 25616 873 25634 907
rect 25564 857 25634 873
rect 25694 907 25764 963
rect 25694 873 25712 907
rect 25746 873 25764 907
rect 25694 857 25764 873
rect 25824 907 25894 963
rect 25824 873 25842 907
rect 25876 873 25894 907
rect 25824 857 25894 873
rect 25954 907 26024 963
rect 25954 873 25972 907
rect 26006 873 26024 907
rect 25954 857 26024 873
rect 26084 907 26154 963
rect 26084 873 26102 907
rect 26136 873 26154 907
rect 26084 857 26154 873
rect 26214 907 26284 963
rect 26214 873 26232 907
rect 26266 873 26284 907
rect 26214 857 26284 873
rect 26344 907 26414 963
rect 26344 873 26362 907
rect 26396 873 26414 907
rect 26344 857 26414 873
rect 26474 907 26544 963
rect 26474 873 26492 907
rect 26526 873 26544 907
rect 26474 857 26544 873
rect 26604 907 26674 963
rect 26604 873 26622 907
rect 26656 873 26674 907
rect 26604 857 26674 873
rect 26734 907 26804 963
rect 26734 873 26752 907
rect 26786 873 26804 907
rect 26734 857 26804 873
rect 26864 907 26934 963
rect 26864 873 26882 907
rect 26916 873 26934 907
rect 26864 857 26934 873
rect 26994 907 27064 963
rect 26994 873 27012 907
rect 27046 873 27064 907
rect 26994 857 27064 873
<< polycont >>
rect 13080 5319 13114 5353
rect 13210 5319 13244 5353
rect 13340 5319 13374 5353
rect 13470 5319 13504 5353
rect 13600 5319 13634 5353
rect 13730 5319 13764 5353
rect 13860 5319 13894 5353
rect 13990 5319 14024 5353
rect 14120 5319 14154 5353
rect 14250 5319 14284 5353
rect 14380 5319 14414 5353
rect 14510 5319 14544 5353
rect 14640 5319 14674 5353
rect 14770 5319 14804 5353
rect 14900 5319 14934 5353
rect 15030 5319 15064 5353
rect 24672 5319 24706 5353
rect 24802 5319 24836 5353
rect 24932 5319 24966 5353
rect 25062 5319 25096 5353
rect 25192 5319 25226 5353
rect 25322 5319 25356 5353
rect 25452 5319 25486 5353
rect 25582 5319 25616 5353
rect 25712 5319 25746 5353
rect 25842 5319 25876 5353
rect 25972 5319 26006 5353
rect 26102 5319 26136 5353
rect 26232 5319 26266 5353
rect 26362 5319 26396 5353
rect 26492 5319 26526 5353
rect 26622 5319 26656 5353
rect 15404 4790 15438 4824
rect 15472 4790 15506 4824
rect 26996 4790 27030 4824
rect 27064 4790 27098 4824
rect 13244 4074 13278 4108
rect 13634 4074 13668 4108
rect 14024 4074 14058 4108
rect 14414 4074 14448 4108
rect 14804 4074 14838 4108
rect 15249 4074 15283 4108
rect 13860 3917 13894 3951
rect 14640 3917 14674 3951
rect 24836 4074 24870 4108
rect 25226 4074 25260 4108
rect 25616 4074 25650 4108
rect 26006 4074 26040 4108
rect 26396 4074 26430 4108
rect 26841 4074 26875 4108
rect 25452 3917 25486 3951
rect 26232 3917 26266 3951
rect 13012 3229 13046 3263
rect 13210 3229 13244 3263
rect 13340 3229 13374 3263
rect 13470 3229 13504 3263
rect 13600 3229 13634 3263
rect 13730 3229 13764 3263
rect 13860 3229 13894 3263
rect 13990 3229 14024 3263
rect 14120 3229 14154 3263
rect 14250 3229 14284 3263
rect 14380 3229 14414 3263
rect 14510 3229 14544 3263
rect 14640 3229 14674 3263
rect 14770 3229 14804 3263
rect 14900 3229 14934 3263
rect 15030 3229 15064 3263
rect 24604 3229 24638 3263
rect 24802 3229 24836 3263
rect 24932 3229 24966 3263
rect 25062 3229 25096 3263
rect 25192 3229 25226 3263
rect 25322 3229 25356 3263
rect 25452 3229 25486 3263
rect 25582 3229 25616 3263
rect 25712 3229 25746 3263
rect 25842 3229 25876 3263
rect 25972 3229 26006 3263
rect 26102 3229 26136 3263
rect 26232 3229 26266 3263
rect 26362 3229 26396 3263
rect 26492 3229 26526 3263
rect 26622 3229 26656 3263
rect 13210 2963 13244 2997
rect 13340 2963 13374 2997
rect 13470 2963 13504 2997
rect 13600 2963 13634 2997
rect 13730 2963 13764 2997
rect 13860 2963 13894 2997
rect 13990 2963 14024 2997
rect 14120 2963 14154 2997
rect 14250 2963 14284 2997
rect 14380 2963 14414 2997
rect 14510 2963 14544 2997
rect 14640 2963 14674 2997
rect 14770 2963 14804 2997
rect 14900 2963 14934 2997
rect 15030 2963 15064 2997
rect 15160 2963 15194 2997
rect 15290 2963 15324 2997
rect 15420 2963 15454 2997
rect 24802 2963 24836 2997
rect 24932 2963 24966 2997
rect 25062 2963 25096 2997
rect 25192 2963 25226 2997
rect 25322 2963 25356 2997
rect 25452 2963 25486 2997
rect 25582 2963 25616 2997
rect 25712 2963 25746 2997
rect 25842 2963 25876 2997
rect 25972 2963 26006 2997
rect 26102 2963 26136 2997
rect 26232 2963 26266 2997
rect 26362 2963 26396 2997
rect 26492 2963 26526 2997
rect 26622 2963 26656 2997
rect 26752 2963 26786 2997
rect 26882 2963 26916 2997
rect 27012 2963 27046 2997
rect 13210 2275 13244 2309
rect 13600 2275 13634 2309
rect 14380 2275 14414 2309
rect 15160 2275 15194 2309
rect 24802 2275 24836 2309
rect 25192 2275 25226 2309
rect 25972 2275 26006 2309
rect 26752 2275 26786 2309
rect 13436 2118 13470 2152
rect 13826 2118 13860 2152
rect 14216 2118 14250 2152
rect 14606 2118 14640 2152
rect 14996 2118 15030 2152
rect 15386 2118 15420 2152
rect 25028 2118 25062 2152
rect 25418 2118 25452 2152
rect 25808 2118 25842 2152
rect 26198 2118 26232 2152
rect 26588 2118 26622 2152
rect 26978 2118 27012 2152
rect 13210 873 13244 907
rect 13340 873 13374 907
rect 13470 873 13504 907
rect 13600 873 13634 907
rect 13730 873 13764 907
rect 13860 873 13894 907
rect 13990 873 14024 907
rect 14120 873 14154 907
rect 14250 873 14284 907
rect 14380 873 14414 907
rect 14510 873 14544 907
rect 14640 873 14674 907
rect 14770 873 14804 907
rect 14900 873 14934 907
rect 15030 873 15064 907
rect 15160 873 15194 907
rect 15290 873 15324 907
rect 15420 873 15454 907
rect 24802 873 24836 907
rect 24932 873 24966 907
rect 25062 873 25096 907
rect 25192 873 25226 907
rect 25322 873 25356 907
rect 25452 873 25486 907
rect 25582 873 25616 907
rect 25712 873 25746 907
rect 25842 873 25876 907
rect 25972 873 26006 907
rect 26102 873 26136 907
rect 26232 873 26266 907
rect 26362 873 26396 907
rect 26492 873 26526 907
rect 26622 873 26656 907
rect 26752 873 26786 907
rect 26882 873 26916 907
rect 27012 873 27046 907
<< locali >>
rect 12998 5486 15112 5509
rect 12998 5452 13022 5486
rect 13056 5452 13104 5486
rect 13138 5452 13196 5486
rect 13238 5452 13268 5486
rect 13306 5452 13340 5486
rect 13374 5452 13408 5486
rect 13446 5452 13476 5486
rect 13518 5452 13586 5486
rect 13628 5452 13658 5486
rect 13696 5452 13730 5486
rect 13764 5452 13798 5486
rect 13836 5452 13866 5486
rect 13908 5452 13976 5486
rect 14018 5452 14048 5486
rect 14086 5452 14120 5486
rect 14154 5452 14188 5486
rect 14226 5452 14256 5486
rect 14298 5452 14366 5486
rect 14408 5452 14438 5486
rect 14476 5452 14510 5486
rect 14544 5452 14578 5486
rect 14616 5452 14646 5486
rect 14688 5452 14756 5486
rect 14798 5452 14828 5486
rect 14866 5452 14900 5486
rect 14934 5452 14968 5486
rect 15006 5452 15036 5486
rect 15078 5452 15112 5486
rect 12998 5429 15112 5452
rect 24590 5486 26704 5509
rect 24590 5452 24614 5486
rect 24648 5452 24696 5486
rect 24730 5452 24788 5486
rect 24830 5452 24860 5486
rect 24898 5452 24932 5486
rect 24966 5452 25000 5486
rect 25038 5452 25068 5486
rect 25110 5452 25178 5486
rect 25220 5452 25250 5486
rect 25288 5452 25322 5486
rect 25356 5452 25390 5486
rect 25428 5452 25458 5486
rect 25500 5452 25568 5486
rect 25610 5452 25640 5486
rect 25678 5452 25712 5486
rect 25746 5452 25780 5486
rect 25818 5452 25848 5486
rect 25890 5452 25958 5486
rect 26000 5452 26030 5486
rect 26068 5452 26102 5486
rect 26136 5452 26170 5486
rect 26208 5452 26238 5486
rect 26280 5452 26348 5486
rect 26390 5452 26420 5486
rect 26458 5452 26492 5486
rect 26526 5452 26560 5486
rect 26598 5452 26628 5486
rect 26670 5452 26704 5486
rect 24590 5429 26704 5452
rect 13064 5319 13080 5353
rect 13114 5319 13130 5353
rect 13194 5319 13210 5353
rect 13244 5319 13260 5353
rect 13324 5319 13340 5353
rect 13374 5319 13390 5353
rect 13454 5319 13470 5353
rect 13504 5319 13520 5353
rect 13584 5319 13600 5353
rect 13634 5319 13650 5353
rect 13714 5319 13730 5353
rect 13764 5319 13780 5353
rect 13844 5319 13860 5353
rect 13894 5319 13910 5353
rect 13974 5319 13990 5353
rect 14024 5319 14040 5353
rect 14104 5319 14120 5353
rect 14154 5319 14170 5353
rect 14234 5319 14250 5353
rect 14284 5319 14300 5353
rect 14364 5319 14380 5353
rect 14414 5319 14430 5353
rect 14494 5319 14510 5353
rect 14544 5319 14560 5353
rect 14624 5319 14640 5353
rect 14674 5319 14690 5353
rect 14754 5319 14770 5353
rect 14804 5319 14820 5353
rect 14884 5319 14900 5353
rect 14934 5319 14950 5353
rect 15014 5319 15030 5353
rect 15064 5319 15080 5353
rect 24656 5319 24672 5353
rect 24706 5319 24722 5353
rect 24786 5319 24802 5353
rect 24836 5319 24852 5353
rect 24916 5319 24932 5353
rect 24966 5319 24982 5353
rect 25046 5319 25062 5353
rect 25096 5319 25112 5353
rect 25176 5319 25192 5353
rect 25226 5319 25242 5353
rect 25306 5319 25322 5353
rect 25356 5319 25372 5353
rect 25436 5319 25452 5353
rect 25486 5319 25502 5353
rect 25566 5319 25582 5353
rect 25616 5319 25632 5353
rect 25696 5319 25712 5353
rect 25746 5319 25762 5353
rect 25826 5319 25842 5353
rect 25876 5319 25892 5353
rect 25956 5319 25972 5353
rect 26006 5319 26022 5353
rect 26086 5319 26102 5353
rect 26136 5319 26152 5353
rect 26216 5319 26232 5353
rect 26266 5319 26282 5353
rect 26346 5319 26362 5353
rect 26396 5319 26412 5353
rect 26476 5319 26492 5353
rect 26526 5319 26542 5353
rect 26606 5319 26622 5353
rect 26656 5319 26672 5353
rect 13015 5224 13049 5240
rect 13015 5152 13049 5190
rect 13015 5080 13049 5118
rect 13015 5008 13049 5046
rect 13015 4936 13049 4974
rect 13015 4886 13049 4902
rect 13145 5224 13179 5240
rect 13145 5152 13179 5190
rect 13145 5080 13179 5118
rect 13145 5008 13179 5046
rect 13145 4936 13179 4974
rect 13145 4886 13179 4902
rect 13275 5224 13309 5240
rect 13275 5152 13309 5190
rect 13275 5080 13309 5118
rect 13275 5008 13309 5046
rect 13275 4936 13309 4974
rect 13275 4886 13309 4902
rect 13405 5224 13439 5240
rect 13405 5152 13439 5190
rect 13405 5080 13439 5118
rect 13405 5008 13439 5046
rect 13405 4936 13439 4974
rect 13405 4886 13439 4902
rect 13535 5224 13569 5240
rect 13535 5152 13569 5190
rect 13535 5080 13569 5118
rect 13535 5008 13569 5046
rect 13535 4936 13569 4974
rect 13535 4886 13569 4902
rect 13665 5224 13699 5240
rect 13665 5152 13699 5190
rect 13665 5080 13699 5118
rect 13665 5008 13699 5046
rect 13665 4936 13699 4974
rect 13665 4886 13699 4902
rect 13795 5224 13829 5240
rect 13795 5152 13829 5190
rect 13795 5080 13829 5118
rect 13795 5008 13829 5046
rect 13795 4936 13829 4974
rect 13795 4886 13829 4902
rect 13925 5224 13959 5240
rect 13925 5152 13959 5190
rect 13925 5080 13959 5118
rect 13925 5008 13959 5046
rect 13925 4936 13959 4974
rect 13925 4886 13959 4902
rect 14055 5224 14089 5240
rect 14055 5152 14089 5190
rect 14055 5080 14089 5118
rect 14055 5008 14089 5046
rect 14055 4936 14089 4974
rect 14055 4886 14089 4902
rect 14185 5224 14219 5240
rect 14185 5152 14219 5190
rect 14185 5080 14219 5118
rect 14185 5008 14219 5046
rect 14185 4936 14219 4974
rect 14185 4886 14219 4902
rect 14315 5224 14349 5240
rect 14315 5152 14349 5190
rect 14315 5080 14349 5118
rect 14315 5008 14349 5046
rect 14315 4936 14349 4974
rect 14315 4886 14349 4902
rect 14445 5224 14479 5240
rect 14445 5152 14479 5190
rect 14445 5080 14479 5118
rect 14445 5008 14479 5046
rect 14445 4936 14479 4974
rect 14445 4886 14479 4902
rect 14575 5224 14609 5240
rect 14575 5152 14609 5190
rect 14575 5080 14609 5118
rect 14575 5008 14609 5046
rect 14575 4936 14609 4974
rect 14575 4886 14609 4902
rect 14705 5224 14739 5240
rect 14705 5152 14739 5190
rect 14705 5080 14739 5118
rect 14705 5008 14739 5046
rect 14705 4936 14739 4974
rect 14705 4886 14739 4902
rect 14835 5224 14869 5240
rect 14835 5152 14869 5190
rect 14835 5080 14869 5118
rect 14835 5008 14869 5046
rect 14835 4936 14869 4974
rect 14835 4886 14869 4902
rect 14965 5224 14999 5240
rect 14965 5152 14999 5190
rect 14965 5080 14999 5118
rect 14965 5008 14999 5046
rect 14965 4936 14999 4974
rect 14965 4886 14999 4902
rect 15095 5224 15129 5240
rect 15095 5152 15129 5190
rect 15095 5080 15129 5118
rect 15095 5008 15129 5046
rect 15095 4936 15129 4974
rect 24607 5224 24641 5240
rect 24607 5152 24641 5190
rect 24607 5080 24641 5118
rect 24607 5008 24641 5046
rect 24607 4936 24641 4974
rect 15095 4886 15129 4902
rect 15284 4915 15524 4927
rect 15284 4881 15315 4915
rect 15353 4881 15387 4915
rect 15421 4881 15455 4915
rect 15493 4881 15524 4915
rect 24607 4886 24641 4902
rect 24737 5224 24771 5240
rect 24737 5152 24771 5190
rect 24737 5080 24771 5118
rect 24737 5008 24771 5046
rect 24737 4936 24771 4974
rect 24737 4886 24771 4902
rect 24867 5224 24901 5240
rect 24867 5152 24901 5190
rect 24867 5080 24901 5118
rect 24867 5008 24901 5046
rect 24867 4936 24901 4974
rect 24867 4886 24901 4902
rect 24997 5224 25031 5240
rect 24997 5152 25031 5190
rect 24997 5080 25031 5118
rect 24997 5008 25031 5046
rect 24997 4936 25031 4974
rect 24997 4886 25031 4902
rect 25127 5224 25161 5240
rect 25127 5152 25161 5190
rect 25127 5080 25161 5118
rect 25127 5008 25161 5046
rect 25127 4936 25161 4974
rect 25127 4886 25161 4902
rect 25257 5224 25291 5240
rect 25257 5152 25291 5190
rect 25257 5080 25291 5118
rect 25257 5008 25291 5046
rect 25257 4936 25291 4974
rect 25257 4886 25291 4902
rect 25387 5224 25421 5240
rect 25387 5152 25421 5190
rect 25387 5080 25421 5118
rect 25387 5008 25421 5046
rect 25387 4936 25421 4974
rect 25387 4886 25421 4902
rect 25517 5224 25551 5240
rect 25517 5152 25551 5190
rect 25517 5080 25551 5118
rect 25517 5008 25551 5046
rect 25517 4936 25551 4974
rect 25517 4886 25551 4902
rect 25647 5224 25681 5240
rect 25647 5152 25681 5190
rect 25647 5080 25681 5118
rect 25647 5008 25681 5046
rect 25647 4936 25681 4974
rect 25647 4886 25681 4902
rect 25777 5224 25811 5240
rect 25777 5152 25811 5190
rect 25777 5080 25811 5118
rect 25777 5008 25811 5046
rect 25777 4936 25811 4974
rect 25777 4886 25811 4902
rect 25907 5224 25941 5240
rect 25907 5152 25941 5190
rect 25907 5080 25941 5118
rect 25907 5008 25941 5046
rect 25907 4936 25941 4974
rect 25907 4886 25941 4902
rect 26037 5224 26071 5240
rect 26037 5152 26071 5190
rect 26037 5080 26071 5118
rect 26037 5008 26071 5046
rect 26037 4936 26071 4974
rect 26037 4886 26071 4902
rect 26167 5224 26201 5240
rect 26167 5152 26201 5190
rect 26167 5080 26201 5118
rect 26167 5008 26201 5046
rect 26167 4936 26201 4974
rect 26167 4886 26201 4902
rect 26297 5224 26331 5240
rect 26297 5152 26331 5190
rect 26297 5080 26331 5118
rect 26297 5008 26331 5046
rect 26297 4936 26331 4974
rect 26297 4886 26331 4902
rect 26427 5224 26461 5240
rect 26427 5152 26461 5190
rect 26427 5080 26461 5118
rect 26427 5008 26461 5046
rect 26427 4936 26461 4974
rect 26427 4886 26461 4902
rect 26557 5224 26591 5240
rect 26557 5152 26591 5190
rect 26557 5080 26591 5118
rect 26557 5008 26591 5046
rect 26557 4936 26591 4974
rect 26557 4886 26591 4902
rect 26687 5224 26721 5240
rect 26687 5152 26721 5190
rect 26687 5080 26721 5118
rect 26687 5008 26721 5046
rect 26687 4936 26721 4974
rect 26687 4886 26721 4902
rect 26876 4915 27116 4927
rect 15284 4869 15524 4881
rect 26876 4881 26907 4915
rect 26945 4881 26979 4915
rect 27013 4881 27047 4915
rect 27085 4881 27116 4915
rect 26876 4869 27116 4881
rect 15375 4824 15535 4834
rect 15375 4790 15402 4824
rect 15438 4790 15472 4824
rect 15508 4790 15535 4824
rect 15375 4780 15535 4790
rect 26967 4824 27127 4834
rect 26967 4790 26994 4824
rect 27030 4790 27064 4824
rect 27100 4790 27127 4824
rect 26967 4780 27127 4790
rect 13275 4676 13309 4692
rect 13275 4604 13309 4642
rect 13275 4532 13309 4570
rect 13275 4460 13309 4498
rect 13275 4388 13309 4426
rect 13275 4338 13309 4354
rect 13405 4676 13439 4692
rect 13405 4604 13439 4642
rect 13405 4532 13439 4570
rect 13405 4460 13439 4498
rect 13405 4388 13439 4426
rect 13405 4338 13439 4354
rect 13665 4676 13699 4692
rect 13665 4604 13699 4642
rect 13665 4532 13699 4570
rect 13665 4460 13699 4498
rect 13665 4388 13699 4426
rect 13665 4338 13699 4354
rect 13795 4676 13829 4692
rect 13795 4604 13829 4642
rect 13795 4532 13829 4570
rect 13795 4460 13829 4498
rect 13795 4388 13829 4426
rect 13795 4338 13829 4354
rect 14055 4676 14089 4692
rect 14055 4604 14089 4642
rect 14055 4532 14089 4570
rect 14055 4460 14089 4498
rect 14055 4388 14089 4426
rect 14055 4338 14089 4354
rect 14185 4676 14219 4692
rect 14185 4604 14219 4642
rect 14185 4532 14219 4570
rect 14185 4460 14219 4498
rect 14185 4388 14219 4426
rect 14185 4338 14219 4354
rect 14445 4676 14479 4692
rect 14445 4604 14479 4642
rect 14445 4532 14479 4570
rect 14445 4460 14479 4498
rect 14445 4388 14479 4426
rect 14445 4338 14479 4354
rect 14575 4676 14609 4692
rect 14575 4604 14609 4642
rect 14575 4532 14609 4570
rect 14575 4460 14609 4498
rect 14575 4388 14609 4426
rect 14575 4338 14609 4354
rect 14835 4676 14869 4692
rect 14835 4604 14869 4642
rect 14835 4532 14869 4570
rect 14835 4460 14869 4498
rect 14835 4388 14869 4426
rect 14835 4338 14869 4354
rect 14965 4676 14999 4692
rect 14965 4604 14999 4642
rect 14965 4532 14999 4570
rect 14965 4460 14999 4498
rect 14965 4388 14999 4426
rect 14965 4338 14999 4354
rect 15209 4676 15243 4692
rect 15209 4604 15243 4642
rect 15209 4532 15243 4570
rect 15209 4460 15243 4498
rect 15209 4388 15243 4426
rect 15209 4338 15243 4354
rect 15299 4676 15333 4692
rect 15299 4604 15333 4642
rect 15299 4532 15333 4570
rect 15299 4460 15333 4498
rect 15299 4388 15333 4426
rect 15299 4338 15333 4354
rect 15389 4676 15423 4692
rect 15389 4604 15423 4642
rect 15389 4532 15423 4570
rect 15389 4460 15423 4498
rect 15389 4388 15423 4426
rect 15389 4338 15423 4354
rect 15479 4676 15513 4692
rect 15479 4604 15513 4642
rect 15479 4532 15513 4570
rect 15479 4460 15513 4498
rect 15479 4388 15513 4426
rect 15479 4338 15513 4354
rect 15569 4676 15603 4692
rect 15569 4604 15603 4642
rect 15569 4532 15603 4570
rect 15569 4460 15603 4498
rect 15569 4388 15603 4426
rect 15569 4338 15603 4354
rect 24867 4676 24901 4692
rect 24867 4604 24901 4642
rect 24867 4532 24901 4570
rect 24867 4460 24901 4498
rect 24867 4388 24901 4426
rect 24867 4338 24901 4354
rect 24997 4676 25031 4692
rect 24997 4604 25031 4642
rect 24997 4532 25031 4570
rect 24997 4460 25031 4498
rect 24997 4388 25031 4426
rect 24997 4338 25031 4354
rect 25257 4676 25291 4692
rect 25257 4604 25291 4642
rect 25257 4532 25291 4570
rect 25257 4460 25291 4498
rect 25257 4388 25291 4426
rect 25257 4338 25291 4354
rect 25387 4676 25421 4692
rect 25387 4604 25421 4642
rect 25387 4532 25421 4570
rect 25387 4460 25421 4498
rect 25387 4388 25421 4426
rect 25387 4338 25421 4354
rect 25647 4676 25681 4692
rect 25647 4604 25681 4642
rect 25647 4532 25681 4570
rect 25647 4460 25681 4498
rect 25647 4388 25681 4426
rect 25647 4338 25681 4354
rect 25777 4676 25811 4692
rect 25777 4604 25811 4642
rect 25777 4532 25811 4570
rect 25777 4460 25811 4498
rect 25777 4388 25811 4426
rect 25777 4338 25811 4354
rect 26037 4676 26071 4692
rect 26037 4604 26071 4642
rect 26037 4532 26071 4570
rect 26037 4460 26071 4498
rect 26037 4388 26071 4426
rect 26037 4338 26071 4354
rect 26167 4676 26201 4692
rect 26167 4604 26201 4642
rect 26167 4532 26201 4570
rect 26167 4460 26201 4498
rect 26167 4388 26201 4426
rect 26167 4338 26201 4354
rect 26427 4676 26461 4692
rect 26427 4604 26461 4642
rect 26427 4532 26461 4570
rect 26427 4460 26461 4498
rect 26427 4388 26461 4426
rect 26427 4338 26461 4354
rect 26557 4676 26591 4692
rect 26557 4604 26591 4642
rect 26557 4532 26591 4570
rect 26557 4460 26591 4498
rect 26557 4388 26591 4426
rect 26557 4338 26591 4354
rect 26801 4676 26835 4692
rect 26801 4604 26835 4642
rect 26801 4532 26835 4570
rect 26801 4460 26835 4498
rect 26801 4388 26835 4426
rect 26801 4338 26835 4354
rect 26891 4676 26925 4692
rect 26891 4604 26925 4642
rect 26891 4532 26925 4570
rect 26891 4460 26925 4498
rect 26891 4388 26925 4426
rect 26891 4338 26925 4354
rect 26981 4676 27015 4692
rect 26981 4604 27015 4642
rect 26981 4532 27015 4570
rect 26981 4460 27015 4498
rect 26981 4388 27015 4426
rect 26981 4338 27015 4354
rect 27071 4676 27105 4692
rect 27071 4604 27105 4642
rect 27071 4532 27105 4570
rect 27071 4460 27105 4498
rect 27071 4388 27105 4426
rect 27071 4338 27105 4354
rect 27161 4676 27195 4692
rect 27161 4604 27195 4642
rect 27161 4532 27195 4570
rect 27161 4460 27195 4498
rect 27161 4388 27195 4426
rect 27161 4338 27195 4354
rect 13228 4108 13294 4123
rect 13228 4074 13244 4108
rect 13278 4074 13294 4108
rect 13228 4059 13294 4074
rect 13618 4108 13684 4123
rect 13618 4074 13634 4108
rect 13668 4074 13684 4108
rect 13618 4059 13684 4074
rect 14008 4108 14074 4123
rect 14008 4074 14024 4108
rect 14058 4074 14074 4108
rect 14008 4059 14074 4074
rect 14398 4108 14464 4123
rect 14398 4074 14414 4108
rect 14448 4074 14464 4108
rect 14398 4059 14464 4074
rect 14788 4108 14854 4123
rect 14788 4074 14804 4108
rect 14838 4074 14854 4108
rect 14788 4059 14854 4074
rect 15233 4108 15299 4118
rect 15233 4074 15249 4108
rect 15283 4074 15299 4108
rect 15233 4064 15299 4074
rect 24820 4108 24886 4123
rect 24820 4074 24836 4108
rect 24870 4074 24886 4108
rect 24820 4059 24886 4074
rect 25210 4108 25276 4123
rect 25210 4074 25226 4108
rect 25260 4074 25276 4108
rect 25210 4059 25276 4074
rect 25600 4108 25666 4123
rect 25600 4074 25616 4108
rect 25650 4074 25666 4108
rect 25600 4059 25666 4074
rect 25990 4108 26056 4123
rect 25990 4074 26006 4108
rect 26040 4074 26056 4108
rect 25990 4059 26056 4074
rect 26380 4108 26446 4123
rect 26380 4074 26396 4108
rect 26430 4074 26446 4108
rect 26380 4059 26446 4074
rect 26825 4108 26891 4118
rect 26825 4074 26841 4108
rect 26875 4074 26891 4108
rect 26825 4064 26891 4074
rect 13842 3951 13912 3961
rect 13842 3917 13860 3951
rect 13894 3917 13912 3951
rect 13842 3907 13912 3917
rect 14622 3951 14692 3961
rect 14622 3917 14640 3951
rect 14674 3917 14692 3951
rect 14622 3907 14692 3917
rect 25434 3951 25504 3961
rect 25434 3917 25452 3951
rect 25486 3917 25504 3951
rect 25434 3907 25504 3917
rect 26214 3951 26284 3961
rect 26214 3917 26232 3951
rect 26266 3917 26284 3951
rect 26214 3907 26284 3917
rect 13275 3820 13309 3836
rect 13275 3748 13309 3786
rect 13275 3698 13309 3714
rect 13405 3820 13439 3836
rect 13405 3748 13439 3786
rect 13405 3698 13439 3714
rect 13535 3820 13569 3836
rect 13535 3748 13569 3786
rect 13535 3698 13569 3714
rect 13665 3820 13699 3836
rect 13665 3748 13699 3786
rect 13665 3698 13699 3714
rect 13795 3820 13829 3836
rect 13795 3748 13829 3786
rect 13795 3698 13829 3714
rect 13925 3820 13959 3836
rect 13925 3748 13959 3786
rect 13925 3698 13959 3714
rect 14055 3820 14089 3836
rect 14055 3748 14089 3786
rect 14055 3698 14089 3714
rect 14185 3820 14219 3836
rect 14185 3748 14219 3786
rect 14185 3698 14219 3714
rect 14315 3820 14349 3836
rect 14315 3748 14349 3786
rect 14315 3698 14349 3714
rect 14445 3820 14479 3836
rect 14445 3748 14479 3786
rect 14445 3698 14479 3714
rect 14575 3820 14609 3836
rect 14575 3748 14609 3786
rect 14575 3698 14609 3714
rect 14705 3820 14739 3836
rect 14705 3748 14739 3786
rect 14705 3698 14739 3714
rect 14835 3820 14869 3836
rect 14835 3748 14869 3786
rect 14835 3698 14869 3714
rect 14965 3820 14999 3836
rect 14965 3748 14999 3786
rect 14965 3698 14999 3714
rect 15095 3820 15129 3836
rect 15095 3748 15129 3786
rect 15095 3698 15129 3714
rect 15209 3820 15243 3836
rect 15209 3748 15243 3786
rect 15209 3698 15243 3714
rect 15299 3820 15333 3836
rect 15299 3748 15333 3786
rect 15299 3698 15333 3714
rect 15389 3820 15423 3836
rect 15389 3748 15423 3786
rect 15389 3698 15423 3714
rect 15479 3820 15513 3836
rect 15479 3748 15513 3786
rect 15479 3698 15513 3714
rect 15569 3820 15603 3836
rect 15569 3748 15603 3786
rect 15569 3698 15603 3714
rect 24867 3820 24901 3836
rect 24867 3748 24901 3786
rect 24867 3698 24901 3714
rect 24997 3820 25031 3836
rect 24997 3748 25031 3786
rect 24997 3698 25031 3714
rect 25127 3820 25161 3836
rect 25127 3748 25161 3786
rect 25127 3698 25161 3714
rect 25257 3820 25291 3836
rect 25257 3748 25291 3786
rect 25257 3698 25291 3714
rect 25387 3820 25421 3836
rect 25387 3748 25421 3786
rect 25387 3698 25421 3714
rect 25517 3820 25551 3836
rect 25517 3748 25551 3786
rect 25517 3698 25551 3714
rect 25647 3820 25681 3836
rect 25647 3748 25681 3786
rect 25647 3698 25681 3714
rect 25777 3820 25811 3836
rect 25777 3748 25811 3786
rect 25777 3698 25811 3714
rect 25907 3820 25941 3836
rect 25907 3748 25941 3786
rect 25907 3698 25941 3714
rect 26037 3820 26071 3836
rect 26037 3748 26071 3786
rect 26037 3698 26071 3714
rect 26167 3820 26201 3836
rect 26167 3748 26201 3786
rect 26167 3698 26201 3714
rect 26297 3820 26331 3836
rect 26297 3748 26331 3786
rect 26297 3698 26331 3714
rect 26427 3820 26461 3836
rect 26427 3748 26461 3786
rect 26427 3698 26461 3714
rect 26557 3820 26591 3836
rect 26557 3748 26591 3786
rect 26557 3698 26591 3714
rect 26687 3820 26721 3836
rect 26687 3748 26721 3786
rect 26687 3698 26721 3714
rect 26801 3820 26835 3836
rect 26801 3748 26835 3786
rect 26801 3698 26835 3714
rect 26891 3820 26925 3836
rect 26891 3748 26925 3786
rect 26891 3698 26925 3714
rect 26981 3820 27015 3836
rect 26981 3748 27015 3786
rect 26981 3698 27015 3714
rect 27071 3820 27105 3836
rect 27071 3748 27105 3786
rect 27071 3698 27105 3714
rect 27161 3820 27195 3836
rect 27161 3748 27195 3786
rect 27161 3698 27195 3714
rect 15287 3579 15527 3591
rect 15287 3545 15318 3579
rect 15356 3545 15390 3579
rect 15424 3545 15458 3579
rect 15496 3545 15527 3579
rect 15287 3533 15527 3545
rect 26879 3579 27119 3591
rect 26879 3545 26910 3579
rect 26948 3545 26982 3579
rect 27016 3545 27050 3579
rect 27088 3545 27119 3579
rect 26879 3533 27119 3545
rect 13015 3472 13049 3488
rect 13015 3400 13049 3438
rect 13015 3350 13049 3366
rect 13145 3472 13179 3488
rect 13145 3400 13179 3438
rect 13145 3350 13179 3366
rect 13275 3472 13309 3488
rect 13275 3400 13309 3438
rect 13275 3350 13309 3366
rect 13405 3472 13439 3488
rect 13405 3400 13439 3438
rect 13405 3350 13439 3366
rect 13535 3472 13569 3488
rect 13535 3400 13569 3438
rect 13535 3350 13569 3366
rect 13665 3472 13699 3488
rect 13665 3400 13699 3438
rect 13665 3350 13699 3366
rect 13795 3472 13829 3488
rect 13795 3400 13829 3438
rect 13795 3350 13829 3366
rect 13925 3472 13959 3488
rect 13925 3400 13959 3438
rect 13925 3350 13959 3366
rect 14055 3472 14089 3488
rect 14055 3400 14089 3438
rect 14055 3350 14089 3366
rect 14185 3472 14219 3488
rect 14185 3400 14219 3438
rect 14185 3350 14219 3366
rect 14315 3472 14349 3488
rect 14315 3400 14349 3438
rect 14315 3350 14349 3366
rect 14445 3472 14479 3488
rect 14445 3400 14479 3438
rect 14445 3350 14479 3366
rect 14575 3472 14609 3488
rect 14575 3400 14609 3438
rect 14575 3350 14609 3366
rect 14705 3472 14739 3488
rect 14705 3400 14739 3438
rect 14705 3350 14739 3366
rect 14835 3472 14869 3488
rect 14835 3400 14869 3438
rect 14835 3350 14869 3366
rect 14965 3472 14999 3488
rect 14965 3400 14999 3438
rect 14965 3350 14999 3366
rect 15095 3472 15129 3488
rect 15095 3400 15129 3438
rect 15095 3350 15129 3366
rect 24607 3472 24641 3488
rect 24607 3400 24641 3438
rect 24607 3350 24641 3366
rect 24737 3472 24771 3488
rect 24737 3400 24771 3438
rect 24737 3350 24771 3366
rect 24867 3472 24901 3488
rect 24867 3400 24901 3438
rect 24867 3350 24901 3366
rect 24997 3472 25031 3488
rect 24997 3400 25031 3438
rect 24997 3350 25031 3366
rect 25127 3472 25161 3488
rect 25127 3400 25161 3438
rect 25127 3350 25161 3366
rect 25257 3472 25291 3488
rect 25257 3400 25291 3438
rect 25257 3350 25291 3366
rect 25387 3472 25421 3488
rect 25387 3400 25421 3438
rect 25387 3350 25421 3366
rect 25517 3472 25551 3488
rect 25517 3400 25551 3438
rect 25517 3350 25551 3366
rect 25647 3472 25681 3488
rect 25647 3400 25681 3438
rect 25647 3350 25681 3366
rect 25777 3472 25811 3488
rect 25777 3400 25811 3438
rect 25777 3350 25811 3366
rect 25907 3472 25941 3488
rect 25907 3400 25941 3438
rect 25907 3350 25941 3366
rect 26037 3472 26071 3488
rect 26037 3400 26071 3438
rect 26037 3350 26071 3366
rect 26167 3472 26201 3488
rect 26167 3400 26201 3438
rect 26167 3350 26201 3366
rect 26297 3472 26331 3488
rect 26297 3400 26331 3438
rect 26297 3350 26331 3366
rect 26427 3472 26461 3488
rect 26427 3400 26461 3438
rect 26427 3350 26461 3366
rect 26557 3472 26591 3488
rect 26557 3400 26591 3438
rect 26557 3350 26591 3366
rect 26687 3472 26721 3488
rect 26687 3400 26721 3438
rect 26687 3350 26721 3366
rect 12996 3263 13062 3279
rect 24588 3263 24654 3279
rect 12996 3229 13012 3263
rect 13046 3229 13062 3263
rect 13194 3229 13210 3263
rect 13244 3229 13260 3263
rect 13324 3229 13340 3263
rect 13374 3229 13390 3263
rect 13454 3229 13470 3263
rect 13504 3229 13520 3263
rect 13584 3229 13600 3263
rect 13634 3229 13650 3263
rect 13714 3229 13730 3263
rect 13764 3229 13780 3263
rect 13844 3229 13860 3263
rect 13894 3229 13910 3263
rect 13974 3229 13990 3263
rect 14024 3229 14040 3263
rect 14104 3229 14120 3263
rect 14154 3229 14170 3263
rect 14234 3229 14250 3263
rect 14284 3229 14300 3263
rect 14364 3229 14380 3263
rect 14414 3229 14430 3263
rect 14494 3229 14510 3263
rect 14544 3229 14560 3263
rect 14624 3229 14640 3263
rect 14674 3229 14690 3263
rect 14754 3229 14770 3263
rect 14804 3229 14820 3263
rect 14884 3229 14900 3263
rect 14934 3229 14950 3263
rect 15014 3229 15030 3263
rect 15064 3229 15080 3263
rect 24588 3229 24604 3263
rect 24638 3229 24654 3263
rect 24786 3229 24802 3263
rect 24836 3229 24852 3263
rect 24916 3229 24932 3263
rect 24966 3229 24982 3263
rect 25046 3229 25062 3263
rect 25096 3229 25112 3263
rect 25176 3229 25192 3263
rect 25226 3229 25242 3263
rect 25306 3229 25322 3263
rect 25356 3229 25372 3263
rect 25436 3229 25452 3263
rect 25486 3229 25502 3263
rect 25566 3229 25582 3263
rect 25616 3229 25632 3263
rect 25696 3229 25712 3263
rect 25746 3229 25762 3263
rect 25826 3229 25842 3263
rect 25876 3229 25892 3263
rect 25956 3229 25972 3263
rect 26006 3229 26022 3263
rect 26086 3229 26102 3263
rect 26136 3229 26152 3263
rect 26216 3229 26232 3263
rect 26266 3229 26282 3263
rect 26346 3229 26362 3263
rect 26396 3229 26412 3263
rect 26476 3229 26492 3263
rect 26526 3229 26542 3263
rect 26606 3229 26622 3263
rect 26656 3229 26672 3263
rect 12996 3213 13062 3229
rect 24588 3213 24654 3229
rect 12998 3130 15502 3153
rect 12998 3096 13022 3130
rect 13056 3096 13104 3130
rect 13138 3096 13196 3130
rect 13238 3096 13268 3130
rect 13306 3096 13340 3130
rect 13374 3096 13408 3130
rect 13446 3096 13476 3130
rect 13518 3096 13586 3130
rect 13628 3096 13658 3130
rect 13696 3096 13730 3130
rect 13764 3096 13798 3130
rect 13836 3096 13866 3130
rect 13908 3096 13976 3130
rect 14018 3096 14048 3130
rect 14086 3096 14120 3130
rect 14154 3096 14188 3130
rect 14226 3096 14256 3130
rect 14298 3096 14366 3130
rect 14408 3096 14438 3130
rect 14476 3096 14510 3130
rect 14544 3096 14578 3130
rect 14616 3096 14646 3130
rect 14688 3096 14756 3130
rect 14798 3096 14828 3130
rect 14866 3096 14900 3130
rect 14934 3096 14968 3130
rect 15006 3096 15036 3130
rect 15078 3096 15146 3130
rect 15188 3096 15218 3130
rect 15256 3096 15290 3130
rect 15324 3096 15358 3130
rect 15396 3096 15426 3130
rect 15468 3096 15502 3130
rect 12998 3073 15502 3096
rect 24590 3130 27094 3153
rect 24590 3096 24614 3130
rect 24648 3096 24696 3130
rect 24730 3096 24788 3130
rect 24830 3096 24860 3130
rect 24898 3096 24932 3130
rect 24966 3096 25000 3130
rect 25038 3096 25068 3130
rect 25110 3096 25178 3130
rect 25220 3096 25250 3130
rect 25288 3096 25322 3130
rect 25356 3096 25390 3130
rect 25428 3096 25458 3130
rect 25500 3096 25568 3130
rect 25610 3096 25640 3130
rect 25678 3096 25712 3130
rect 25746 3096 25780 3130
rect 25818 3096 25848 3130
rect 25890 3096 25958 3130
rect 26000 3096 26030 3130
rect 26068 3096 26102 3130
rect 26136 3096 26170 3130
rect 26208 3096 26238 3130
rect 26280 3096 26348 3130
rect 26390 3096 26420 3130
rect 26458 3096 26492 3130
rect 26526 3096 26560 3130
rect 26598 3096 26628 3130
rect 26670 3096 26738 3130
rect 26780 3096 26810 3130
rect 26848 3096 26882 3130
rect 26916 3096 26950 3130
rect 26988 3096 27018 3130
rect 27060 3096 27094 3130
rect 24590 3073 27094 3096
rect 13194 2963 13210 2997
rect 13244 2963 13260 2997
rect 13324 2963 13340 2997
rect 13374 2963 13390 2997
rect 13454 2963 13470 2997
rect 13504 2963 13520 2997
rect 13584 2963 13600 2997
rect 13634 2963 13650 2997
rect 13714 2963 13730 2997
rect 13764 2963 13780 2997
rect 13844 2963 13860 2997
rect 13894 2963 13910 2997
rect 13974 2963 13990 2997
rect 14024 2963 14040 2997
rect 14104 2963 14120 2997
rect 14154 2963 14170 2997
rect 14234 2963 14250 2997
rect 14284 2963 14300 2997
rect 14364 2963 14380 2997
rect 14414 2963 14430 2997
rect 14494 2963 14510 2997
rect 14544 2963 14560 2997
rect 14624 2963 14640 2997
rect 14674 2963 14690 2997
rect 14754 2963 14770 2997
rect 14804 2963 14820 2997
rect 14884 2963 14900 2997
rect 14934 2963 14950 2997
rect 15014 2963 15030 2997
rect 15064 2963 15080 2997
rect 15144 2963 15160 2997
rect 15194 2963 15210 2997
rect 15274 2963 15290 2997
rect 15324 2963 15340 2997
rect 15404 2963 15420 2997
rect 15454 2963 15470 2997
rect 24786 2963 24802 2997
rect 24836 2963 24852 2997
rect 24916 2963 24932 2997
rect 24966 2963 24982 2997
rect 25046 2963 25062 2997
rect 25096 2963 25112 2997
rect 25176 2963 25192 2997
rect 25226 2963 25242 2997
rect 25306 2963 25322 2997
rect 25356 2963 25372 2997
rect 25436 2963 25452 2997
rect 25486 2963 25502 2997
rect 25566 2963 25582 2997
rect 25616 2963 25632 2997
rect 25696 2963 25712 2997
rect 25746 2963 25762 2997
rect 25826 2963 25842 2997
rect 25876 2963 25892 2997
rect 25956 2963 25972 2997
rect 26006 2963 26022 2997
rect 26086 2963 26102 2997
rect 26136 2963 26152 2997
rect 26216 2963 26232 2997
rect 26266 2963 26282 2997
rect 26346 2963 26362 2997
rect 26396 2963 26412 2997
rect 26476 2963 26492 2997
rect 26526 2963 26542 2997
rect 26606 2963 26622 2997
rect 26656 2963 26672 2997
rect 26736 2963 26752 2997
rect 26786 2963 26802 2997
rect 26866 2963 26882 2997
rect 26916 2963 26932 2997
rect 26996 2963 27012 2997
rect 27046 2963 27062 2997
rect 13145 2860 13179 2876
rect 13145 2788 13179 2826
rect 13145 2738 13179 2754
rect 13275 2860 13309 2876
rect 13275 2788 13309 2826
rect 13275 2738 13309 2754
rect 13405 2860 13439 2876
rect 13405 2788 13439 2826
rect 13405 2738 13439 2754
rect 13535 2860 13569 2876
rect 13535 2788 13569 2826
rect 13535 2738 13569 2754
rect 13665 2860 13699 2876
rect 13665 2788 13699 2826
rect 13665 2738 13699 2754
rect 13795 2860 13829 2876
rect 13795 2788 13829 2826
rect 13795 2738 13829 2754
rect 13925 2860 13959 2876
rect 13925 2788 13959 2826
rect 13925 2738 13959 2754
rect 14055 2860 14089 2876
rect 14055 2788 14089 2826
rect 14055 2738 14089 2754
rect 14185 2860 14219 2876
rect 14185 2788 14219 2826
rect 14185 2738 14219 2754
rect 14315 2860 14349 2876
rect 14315 2788 14349 2826
rect 14315 2738 14349 2754
rect 14445 2860 14479 2876
rect 14445 2788 14479 2826
rect 14445 2738 14479 2754
rect 14575 2860 14609 2876
rect 14575 2788 14609 2826
rect 14575 2738 14609 2754
rect 14705 2860 14739 2876
rect 14705 2788 14739 2826
rect 14705 2738 14739 2754
rect 14835 2860 14869 2876
rect 14835 2788 14869 2826
rect 14835 2738 14869 2754
rect 14965 2860 14999 2876
rect 14965 2788 14999 2826
rect 14965 2738 14999 2754
rect 15095 2860 15129 2876
rect 15095 2788 15129 2826
rect 15095 2738 15129 2754
rect 15225 2860 15259 2876
rect 15225 2788 15259 2826
rect 15225 2738 15259 2754
rect 15355 2860 15389 2876
rect 15355 2788 15389 2826
rect 15355 2738 15389 2754
rect 15485 2860 15519 2876
rect 15485 2788 15519 2826
rect 15485 2738 15519 2754
rect 24737 2860 24771 2876
rect 24737 2788 24771 2826
rect 24737 2738 24771 2754
rect 24867 2860 24901 2876
rect 24867 2788 24901 2826
rect 24867 2738 24901 2754
rect 24997 2860 25031 2876
rect 24997 2788 25031 2826
rect 24997 2738 25031 2754
rect 25127 2860 25161 2876
rect 25127 2788 25161 2826
rect 25127 2738 25161 2754
rect 25257 2860 25291 2876
rect 25257 2788 25291 2826
rect 25257 2738 25291 2754
rect 25387 2860 25421 2876
rect 25387 2788 25421 2826
rect 25387 2738 25421 2754
rect 25517 2860 25551 2876
rect 25517 2788 25551 2826
rect 25517 2738 25551 2754
rect 25647 2860 25681 2876
rect 25647 2788 25681 2826
rect 25647 2738 25681 2754
rect 25777 2860 25811 2876
rect 25777 2788 25811 2826
rect 25777 2738 25811 2754
rect 25907 2860 25941 2876
rect 25907 2788 25941 2826
rect 25907 2738 25941 2754
rect 26037 2860 26071 2876
rect 26037 2788 26071 2826
rect 26037 2738 26071 2754
rect 26167 2860 26201 2876
rect 26167 2788 26201 2826
rect 26167 2738 26201 2754
rect 26297 2860 26331 2876
rect 26297 2788 26331 2826
rect 26297 2738 26331 2754
rect 26427 2860 26461 2876
rect 26427 2788 26461 2826
rect 26427 2738 26461 2754
rect 26557 2860 26591 2876
rect 26557 2788 26591 2826
rect 26557 2738 26591 2754
rect 26687 2860 26721 2876
rect 26687 2788 26721 2826
rect 26687 2738 26721 2754
rect 26817 2860 26851 2876
rect 26817 2788 26851 2826
rect 26817 2738 26851 2754
rect 26947 2860 26981 2876
rect 26947 2788 26981 2826
rect 26947 2738 26981 2754
rect 27077 2860 27111 2876
rect 27077 2788 27111 2826
rect 27077 2738 27111 2754
rect 13145 2512 13179 2528
rect 13145 2440 13179 2478
rect 13145 2390 13179 2406
rect 13275 2512 13309 2528
rect 13275 2440 13309 2478
rect 13275 2390 13309 2406
rect 13405 2512 13439 2528
rect 13405 2440 13439 2478
rect 13405 2390 13439 2406
rect 13535 2512 13569 2528
rect 13535 2440 13569 2478
rect 13535 2390 13569 2406
rect 13665 2512 13699 2528
rect 13665 2440 13699 2478
rect 13665 2390 13699 2406
rect 13795 2512 13829 2528
rect 13795 2440 13829 2478
rect 13795 2390 13829 2406
rect 13925 2512 13959 2528
rect 13925 2440 13959 2478
rect 13925 2390 13959 2406
rect 14055 2512 14089 2528
rect 14055 2440 14089 2478
rect 14055 2390 14089 2406
rect 14185 2512 14219 2528
rect 14185 2440 14219 2478
rect 14185 2390 14219 2406
rect 14315 2512 14349 2528
rect 14315 2440 14349 2478
rect 14315 2390 14349 2406
rect 14445 2512 14479 2528
rect 14445 2440 14479 2478
rect 14445 2390 14479 2406
rect 14575 2512 14609 2528
rect 14575 2440 14609 2478
rect 14575 2390 14609 2406
rect 14705 2512 14739 2528
rect 14705 2440 14739 2478
rect 14705 2390 14739 2406
rect 14835 2512 14869 2528
rect 14835 2440 14869 2478
rect 14835 2390 14869 2406
rect 14965 2512 14999 2528
rect 14965 2440 14999 2478
rect 14965 2390 14999 2406
rect 15095 2512 15129 2528
rect 15095 2440 15129 2478
rect 15095 2390 15129 2406
rect 15225 2512 15259 2528
rect 15225 2440 15259 2478
rect 15225 2390 15259 2406
rect 15355 2512 15389 2528
rect 15355 2440 15389 2478
rect 15355 2390 15389 2406
rect 24737 2512 24771 2528
rect 24737 2440 24771 2478
rect 24737 2390 24771 2406
rect 24867 2512 24901 2528
rect 24867 2440 24901 2478
rect 24867 2390 24901 2406
rect 24997 2512 25031 2528
rect 24997 2440 25031 2478
rect 24997 2390 25031 2406
rect 25127 2512 25161 2528
rect 25127 2440 25161 2478
rect 25127 2390 25161 2406
rect 25257 2512 25291 2528
rect 25257 2440 25291 2478
rect 25257 2390 25291 2406
rect 25387 2512 25421 2528
rect 25387 2440 25421 2478
rect 25387 2390 25421 2406
rect 25517 2512 25551 2528
rect 25517 2440 25551 2478
rect 25517 2390 25551 2406
rect 25647 2512 25681 2528
rect 25647 2440 25681 2478
rect 25647 2390 25681 2406
rect 25777 2512 25811 2528
rect 25777 2440 25811 2478
rect 25777 2390 25811 2406
rect 25907 2512 25941 2528
rect 25907 2440 25941 2478
rect 25907 2390 25941 2406
rect 26037 2512 26071 2528
rect 26037 2440 26071 2478
rect 26037 2390 26071 2406
rect 26167 2512 26201 2528
rect 26167 2440 26201 2478
rect 26167 2390 26201 2406
rect 26297 2512 26331 2528
rect 26297 2440 26331 2478
rect 26297 2390 26331 2406
rect 26427 2512 26461 2528
rect 26427 2440 26461 2478
rect 26427 2390 26461 2406
rect 26557 2512 26591 2528
rect 26557 2440 26591 2478
rect 26557 2390 26591 2406
rect 26687 2512 26721 2528
rect 26687 2440 26721 2478
rect 26687 2390 26721 2406
rect 26817 2512 26851 2528
rect 26817 2440 26851 2478
rect 26817 2390 26851 2406
rect 26947 2512 26981 2528
rect 26947 2440 26981 2478
rect 26947 2390 26981 2406
rect 13192 2309 13262 2319
rect 13192 2275 13210 2309
rect 13244 2275 13262 2309
rect 13192 2265 13262 2275
rect 13582 2309 13652 2319
rect 13582 2275 13600 2309
rect 13634 2275 13652 2309
rect 13582 2265 13652 2275
rect 14362 2309 14432 2319
rect 14362 2275 14380 2309
rect 14414 2275 14432 2309
rect 14362 2265 14432 2275
rect 15142 2309 15212 2319
rect 15142 2275 15160 2309
rect 15194 2275 15212 2309
rect 15142 2265 15212 2275
rect 24784 2309 24854 2319
rect 24784 2275 24802 2309
rect 24836 2275 24854 2309
rect 24784 2265 24854 2275
rect 25174 2309 25244 2319
rect 25174 2275 25192 2309
rect 25226 2275 25244 2309
rect 25174 2265 25244 2275
rect 25954 2309 26024 2319
rect 25954 2275 25972 2309
rect 26006 2275 26024 2309
rect 25954 2265 26024 2275
rect 26734 2309 26804 2319
rect 26734 2275 26752 2309
rect 26786 2275 26804 2309
rect 26734 2265 26804 2275
rect 13420 2152 13486 2167
rect 13420 2118 13436 2152
rect 13470 2118 13486 2152
rect 13420 2103 13486 2118
rect 13810 2152 13876 2167
rect 13810 2118 13826 2152
rect 13860 2118 13876 2152
rect 13810 2103 13876 2118
rect 14200 2152 14266 2167
rect 14200 2118 14216 2152
rect 14250 2118 14266 2152
rect 14200 2103 14266 2118
rect 14590 2152 14656 2167
rect 14590 2118 14606 2152
rect 14640 2118 14656 2152
rect 14590 2103 14656 2118
rect 14980 2152 15046 2167
rect 14980 2118 14996 2152
rect 15030 2118 15046 2152
rect 14980 2103 15046 2118
rect 15370 2152 15436 2167
rect 15370 2118 15386 2152
rect 15420 2118 15436 2152
rect 15370 2103 15436 2118
rect 25012 2152 25078 2167
rect 25012 2118 25028 2152
rect 25062 2118 25078 2152
rect 25012 2103 25078 2118
rect 25402 2152 25468 2167
rect 25402 2118 25418 2152
rect 25452 2118 25468 2152
rect 25402 2103 25468 2118
rect 25792 2152 25858 2167
rect 25792 2118 25808 2152
rect 25842 2118 25858 2152
rect 25792 2103 25858 2118
rect 26182 2152 26248 2167
rect 26182 2118 26198 2152
rect 26232 2118 26248 2152
rect 26182 2103 26248 2118
rect 26572 2152 26638 2167
rect 26572 2118 26588 2152
rect 26622 2118 26638 2152
rect 26572 2103 26638 2118
rect 26962 2152 27028 2167
rect 26962 2118 26978 2152
rect 27012 2118 27028 2152
rect 26962 2103 27028 2118
rect 13275 1872 13309 1888
rect 13275 1800 13309 1838
rect 13275 1728 13309 1766
rect 13275 1656 13309 1694
rect 13275 1584 13309 1622
rect 13275 1534 13309 1550
rect 13405 1872 13439 1888
rect 13405 1800 13439 1838
rect 13405 1728 13439 1766
rect 13405 1656 13439 1694
rect 13405 1584 13439 1622
rect 13405 1534 13439 1550
rect 13665 1872 13699 1888
rect 13665 1800 13699 1838
rect 13665 1728 13699 1766
rect 13665 1656 13699 1694
rect 13665 1584 13699 1622
rect 13665 1534 13699 1550
rect 13795 1872 13829 1888
rect 13795 1800 13829 1838
rect 13795 1728 13829 1766
rect 13795 1656 13829 1694
rect 13795 1584 13829 1622
rect 13795 1534 13829 1550
rect 14055 1872 14089 1888
rect 14055 1800 14089 1838
rect 14055 1728 14089 1766
rect 14055 1656 14089 1694
rect 14055 1584 14089 1622
rect 14055 1534 14089 1550
rect 14185 1872 14219 1888
rect 14185 1800 14219 1838
rect 14185 1728 14219 1766
rect 14185 1656 14219 1694
rect 14185 1584 14219 1622
rect 14185 1534 14219 1550
rect 14445 1872 14479 1888
rect 14445 1800 14479 1838
rect 14445 1728 14479 1766
rect 14445 1656 14479 1694
rect 14445 1584 14479 1622
rect 14445 1534 14479 1550
rect 14575 1872 14609 1888
rect 14575 1800 14609 1838
rect 14575 1728 14609 1766
rect 14575 1656 14609 1694
rect 14575 1584 14609 1622
rect 14575 1534 14609 1550
rect 14835 1872 14869 1888
rect 14835 1800 14869 1838
rect 14835 1728 14869 1766
rect 14835 1656 14869 1694
rect 14835 1584 14869 1622
rect 14835 1534 14869 1550
rect 14965 1872 14999 1888
rect 14965 1800 14999 1838
rect 14965 1728 14999 1766
rect 14965 1656 14999 1694
rect 14965 1584 14999 1622
rect 14965 1534 14999 1550
rect 15225 1872 15259 1888
rect 15225 1800 15259 1838
rect 15225 1728 15259 1766
rect 15225 1656 15259 1694
rect 15225 1584 15259 1622
rect 15225 1534 15259 1550
rect 15355 1872 15389 1888
rect 15355 1800 15389 1838
rect 15355 1728 15389 1766
rect 15355 1656 15389 1694
rect 15355 1584 15389 1622
rect 15355 1534 15389 1550
rect 24867 1872 24901 1888
rect 24867 1800 24901 1838
rect 24867 1728 24901 1766
rect 24867 1656 24901 1694
rect 24867 1584 24901 1622
rect 24867 1534 24901 1550
rect 24997 1872 25031 1888
rect 24997 1800 25031 1838
rect 24997 1728 25031 1766
rect 24997 1656 25031 1694
rect 24997 1584 25031 1622
rect 24997 1534 25031 1550
rect 25257 1872 25291 1888
rect 25257 1800 25291 1838
rect 25257 1728 25291 1766
rect 25257 1656 25291 1694
rect 25257 1584 25291 1622
rect 25257 1534 25291 1550
rect 25387 1872 25421 1888
rect 25387 1800 25421 1838
rect 25387 1728 25421 1766
rect 25387 1656 25421 1694
rect 25387 1584 25421 1622
rect 25387 1534 25421 1550
rect 25647 1872 25681 1888
rect 25647 1800 25681 1838
rect 25647 1728 25681 1766
rect 25647 1656 25681 1694
rect 25647 1584 25681 1622
rect 25647 1534 25681 1550
rect 25777 1872 25811 1888
rect 25777 1800 25811 1838
rect 25777 1728 25811 1766
rect 25777 1656 25811 1694
rect 25777 1584 25811 1622
rect 25777 1534 25811 1550
rect 26037 1872 26071 1888
rect 26037 1800 26071 1838
rect 26037 1728 26071 1766
rect 26037 1656 26071 1694
rect 26037 1584 26071 1622
rect 26037 1534 26071 1550
rect 26167 1872 26201 1888
rect 26167 1800 26201 1838
rect 26167 1728 26201 1766
rect 26167 1656 26201 1694
rect 26167 1584 26201 1622
rect 26167 1534 26201 1550
rect 26427 1872 26461 1888
rect 26427 1800 26461 1838
rect 26427 1728 26461 1766
rect 26427 1656 26461 1694
rect 26427 1584 26461 1622
rect 26427 1534 26461 1550
rect 26557 1872 26591 1888
rect 26557 1800 26591 1838
rect 26557 1728 26591 1766
rect 26557 1656 26591 1694
rect 26557 1584 26591 1622
rect 26557 1534 26591 1550
rect 26817 1872 26851 1888
rect 26817 1800 26851 1838
rect 26817 1728 26851 1766
rect 26817 1656 26851 1694
rect 26817 1584 26851 1622
rect 26817 1534 26851 1550
rect 26947 1872 26981 1888
rect 26947 1800 26981 1838
rect 26947 1728 26981 1766
rect 26947 1656 26981 1694
rect 26947 1584 26981 1622
rect 26947 1534 26981 1550
rect 13145 1324 13179 1340
rect 13145 1252 13179 1290
rect 13145 1180 13179 1218
rect 13145 1108 13179 1146
rect 13145 1036 13179 1074
rect 13145 986 13179 1002
rect 13275 1324 13309 1340
rect 13275 1252 13309 1290
rect 13275 1180 13309 1218
rect 13275 1108 13309 1146
rect 13275 1036 13309 1074
rect 13275 986 13309 1002
rect 13405 1324 13439 1340
rect 13405 1252 13439 1290
rect 13405 1180 13439 1218
rect 13405 1108 13439 1146
rect 13405 1036 13439 1074
rect 13405 986 13439 1002
rect 13535 1324 13569 1340
rect 13535 1252 13569 1290
rect 13535 1180 13569 1218
rect 13535 1108 13569 1146
rect 13535 1036 13569 1074
rect 13535 986 13569 1002
rect 13665 1324 13699 1340
rect 13665 1252 13699 1290
rect 13665 1180 13699 1218
rect 13665 1108 13699 1146
rect 13665 1036 13699 1074
rect 13665 986 13699 1002
rect 13795 1324 13829 1340
rect 13795 1252 13829 1290
rect 13795 1180 13829 1218
rect 13795 1108 13829 1146
rect 13795 1036 13829 1074
rect 13795 986 13829 1002
rect 13925 1324 13959 1340
rect 13925 1252 13959 1290
rect 13925 1180 13959 1218
rect 13925 1108 13959 1146
rect 13925 1036 13959 1074
rect 13925 986 13959 1002
rect 14055 1324 14089 1340
rect 14055 1252 14089 1290
rect 14055 1180 14089 1218
rect 14055 1108 14089 1146
rect 14055 1036 14089 1074
rect 14055 986 14089 1002
rect 14185 1324 14219 1340
rect 14185 1252 14219 1290
rect 14185 1180 14219 1218
rect 14185 1108 14219 1146
rect 14185 1036 14219 1074
rect 14185 986 14219 1002
rect 14315 1324 14349 1340
rect 14315 1252 14349 1290
rect 14315 1180 14349 1218
rect 14315 1108 14349 1146
rect 14315 1036 14349 1074
rect 14315 986 14349 1002
rect 14445 1324 14479 1340
rect 14445 1252 14479 1290
rect 14445 1180 14479 1218
rect 14445 1108 14479 1146
rect 14445 1036 14479 1074
rect 14445 986 14479 1002
rect 14575 1324 14609 1340
rect 14575 1252 14609 1290
rect 14575 1180 14609 1218
rect 14575 1108 14609 1146
rect 14575 1036 14609 1074
rect 14575 986 14609 1002
rect 14705 1324 14739 1340
rect 14705 1252 14739 1290
rect 14705 1180 14739 1218
rect 14705 1108 14739 1146
rect 14705 1036 14739 1074
rect 14705 986 14739 1002
rect 14835 1324 14869 1340
rect 14835 1252 14869 1290
rect 14835 1180 14869 1218
rect 14835 1108 14869 1146
rect 14835 1036 14869 1074
rect 14835 986 14869 1002
rect 14965 1324 14999 1340
rect 14965 1252 14999 1290
rect 14965 1180 14999 1218
rect 14965 1108 14999 1146
rect 14965 1036 14999 1074
rect 14965 986 14999 1002
rect 15095 1324 15129 1340
rect 15095 1252 15129 1290
rect 15095 1180 15129 1218
rect 15095 1108 15129 1146
rect 15095 1036 15129 1074
rect 15095 986 15129 1002
rect 15225 1324 15259 1340
rect 15225 1252 15259 1290
rect 15225 1180 15259 1218
rect 15225 1108 15259 1146
rect 15225 1036 15259 1074
rect 15225 986 15259 1002
rect 15355 1324 15389 1340
rect 15355 1252 15389 1290
rect 15355 1180 15389 1218
rect 15355 1108 15389 1146
rect 15355 1036 15389 1074
rect 15355 986 15389 1002
rect 15485 1324 15519 1340
rect 15485 1252 15519 1290
rect 15485 1180 15519 1218
rect 15485 1108 15519 1146
rect 15485 1036 15519 1074
rect 15485 986 15519 1002
rect 24737 1324 24771 1340
rect 24737 1252 24771 1290
rect 24737 1180 24771 1218
rect 24737 1108 24771 1146
rect 24737 1036 24771 1074
rect 24737 986 24771 1002
rect 24867 1324 24901 1340
rect 24867 1252 24901 1290
rect 24867 1180 24901 1218
rect 24867 1108 24901 1146
rect 24867 1036 24901 1074
rect 24867 986 24901 1002
rect 24997 1324 25031 1340
rect 24997 1252 25031 1290
rect 24997 1180 25031 1218
rect 24997 1108 25031 1146
rect 24997 1036 25031 1074
rect 24997 986 25031 1002
rect 25127 1324 25161 1340
rect 25127 1252 25161 1290
rect 25127 1180 25161 1218
rect 25127 1108 25161 1146
rect 25127 1036 25161 1074
rect 25127 986 25161 1002
rect 25257 1324 25291 1340
rect 25257 1252 25291 1290
rect 25257 1180 25291 1218
rect 25257 1108 25291 1146
rect 25257 1036 25291 1074
rect 25257 986 25291 1002
rect 25387 1324 25421 1340
rect 25387 1252 25421 1290
rect 25387 1180 25421 1218
rect 25387 1108 25421 1146
rect 25387 1036 25421 1074
rect 25387 986 25421 1002
rect 25517 1324 25551 1340
rect 25517 1252 25551 1290
rect 25517 1180 25551 1218
rect 25517 1108 25551 1146
rect 25517 1036 25551 1074
rect 25517 986 25551 1002
rect 25647 1324 25681 1340
rect 25647 1252 25681 1290
rect 25647 1180 25681 1218
rect 25647 1108 25681 1146
rect 25647 1036 25681 1074
rect 25647 986 25681 1002
rect 25777 1324 25811 1340
rect 25777 1252 25811 1290
rect 25777 1180 25811 1218
rect 25777 1108 25811 1146
rect 25777 1036 25811 1074
rect 25777 986 25811 1002
rect 25907 1324 25941 1340
rect 25907 1252 25941 1290
rect 25907 1180 25941 1218
rect 25907 1108 25941 1146
rect 25907 1036 25941 1074
rect 25907 986 25941 1002
rect 26037 1324 26071 1340
rect 26037 1252 26071 1290
rect 26037 1180 26071 1218
rect 26037 1108 26071 1146
rect 26037 1036 26071 1074
rect 26037 986 26071 1002
rect 26167 1324 26201 1340
rect 26167 1252 26201 1290
rect 26167 1180 26201 1218
rect 26167 1108 26201 1146
rect 26167 1036 26201 1074
rect 26167 986 26201 1002
rect 26297 1324 26331 1340
rect 26297 1252 26331 1290
rect 26297 1180 26331 1218
rect 26297 1108 26331 1146
rect 26297 1036 26331 1074
rect 26297 986 26331 1002
rect 26427 1324 26461 1340
rect 26427 1252 26461 1290
rect 26427 1180 26461 1218
rect 26427 1108 26461 1146
rect 26427 1036 26461 1074
rect 26427 986 26461 1002
rect 26557 1324 26591 1340
rect 26557 1252 26591 1290
rect 26557 1180 26591 1218
rect 26557 1108 26591 1146
rect 26557 1036 26591 1074
rect 26557 986 26591 1002
rect 26687 1324 26721 1340
rect 26687 1252 26721 1290
rect 26687 1180 26721 1218
rect 26687 1108 26721 1146
rect 26687 1036 26721 1074
rect 26687 986 26721 1002
rect 26817 1324 26851 1340
rect 26817 1252 26851 1290
rect 26817 1180 26851 1218
rect 26817 1108 26851 1146
rect 26817 1036 26851 1074
rect 26817 986 26851 1002
rect 26947 1324 26981 1340
rect 26947 1252 26981 1290
rect 26947 1180 26981 1218
rect 26947 1108 26981 1146
rect 26947 1036 26981 1074
rect 26947 986 26981 1002
rect 27077 1324 27111 1340
rect 27077 1252 27111 1290
rect 27077 1180 27111 1218
rect 27077 1108 27111 1146
rect 27077 1036 27111 1074
rect 27077 986 27111 1002
rect 13194 873 13210 907
rect 13244 873 13260 907
rect 13324 873 13340 907
rect 13374 873 13390 907
rect 13454 873 13470 907
rect 13504 873 13520 907
rect 13584 873 13600 907
rect 13634 873 13650 907
rect 13714 873 13730 907
rect 13764 873 13780 907
rect 13844 873 13860 907
rect 13894 873 13910 907
rect 13974 873 13990 907
rect 14024 873 14040 907
rect 14104 873 14120 907
rect 14154 873 14170 907
rect 14234 873 14250 907
rect 14284 873 14300 907
rect 14364 873 14380 907
rect 14414 873 14430 907
rect 14494 873 14510 907
rect 14544 873 14560 907
rect 14624 873 14640 907
rect 14674 873 14690 907
rect 14754 873 14770 907
rect 14804 873 14820 907
rect 14884 873 14900 907
rect 14934 873 14950 907
rect 15014 873 15030 907
rect 15064 873 15080 907
rect 15144 873 15160 907
rect 15194 873 15210 907
rect 15274 873 15290 907
rect 15324 873 15340 907
rect 15404 873 15420 907
rect 15454 873 15470 907
rect 24786 873 24802 907
rect 24836 873 24852 907
rect 24916 873 24932 907
rect 24966 873 24982 907
rect 25046 873 25062 907
rect 25096 873 25112 907
rect 25176 873 25192 907
rect 25226 873 25242 907
rect 25306 873 25322 907
rect 25356 873 25372 907
rect 25436 873 25452 907
rect 25486 873 25502 907
rect 25566 873 25582 907
rect 25616 873 25632 907
rect 25696 873 25712 907
rect 25746 873 25762 907
rect 25826 873 25842 907
rect 25876 873 25892 907
rect 25956 873 25972 907
rect 26006 873 26022 907
rect 26086 873 26102 907
rect 26136 873 26152 907
rect 26216 873 26232 907
rect 26266 873 26282 907
rect 26346 873 26362 907
rect 26396 873 26412 907
rect 26476 873 26492 907
rect 26526 873 26542 907
rect 26606 873 26622 907
rect 26656 873 26672 907
rect 26736 873 26752 907
rect 26786 873 26802 907
rect 26866 873 26882 907
rect 26916 873 26932 907
rect 26996 873 27012 907
rect 27046 873 27062 907
rect 13162 774 15502 797
rect 13162 740 13196 774
rect 13238 740 13268 774
rect 13306 740 13340 774
rect 13374 740 13408 774
rect 13446 740 13476 774
rect 13518 740 13586 774
rect 13628 740 13658 774
rect 13696 740 13730 774
rect 13764 740 13798 774
rect 13836 740 13866 774
rect 13908 740 13976 774
rect 14018 740 14048 774
rect 14086 740 14120 774
rect 14154 740 14188 774
rect 14226 740 14256 774
rect 14298 740 14366 774
rect 14408 740 14438 774
rect 14476 740 14510 774
rect 14544 740 14578 774
rect 14616 740 14646 774
rect 14688 740 14756 774
rect 14798 740 14828 774
rect 14866 740 14900 774
rect 14934 740 14968 774
rect 15006 740 15036 774
rect 15078 740 15146 774
rect 15188 740 15218 774
rect 15256 740 15290 774
rect 15324 740 15358 774
rect 15396 740 15426 774
rect 15468 740 15502 774
rect 13162 717 15502 740
rect 24754 774 27094 797
rect 24754 740 24788 774
rect 24830 740 24860 774
rect 24898 740 24932 774
rect 24966 740 25000 774
rect 25038 740 25068 774
rect 25110 740 25178 774
rect 25220 740 25250 774
rect 25288 740 25322 774
rect 25356 740 25390 774
rect 25428 740 25458 774
rect 25500 740 25568 774
rect 25610 740 25640 774
rect 25678 740 25712 774
rect 25746 740 25780 774
rect 25818 740 25848 774
rect 25890 740 25958 774
rect 26000 740 26030 774
rect 26068 740 26102 774
rect 26136 740 26170 774
rect 26208 740 26238 774
rect 26280 740 26348 774
rect 26390 740 26420 774
rect 26458 740 26492 774
rect 26526 740 26560 774
rect 26598 740 26628 774
rect 26670 740 26738 774
rect 26780 740 26810 774
rect 26848 740 26882 774
rect 26916 740 26950 774
rect 26988 740 27018 774
rect 27060 740 27094 774
rect 24754 717 27094 740
<< viali >>
rect 13022 5452 13056 5486
rect 13104 5452 13138 5486
rect 13196 5452 13204 5486
rect 13204 5452 13230 5486
rect 13268 5452 13272 5486
rect 13272 5452 13302 5486
rect 13340 5452 13374 5486
rect 13412 5452 13442 5486
rect 13442 5452 13446 5486
rect 13484 5452 13510 5486
rect 13510 5452 13518 5486
rect 13586 5452 13594 5486
rect 13594 5452 13620 5486
rect 13658 5452 13662 5486
rect 13662 5452 13692 5486
rect 13730 5452 13764 5486
rect 13802 5452 13832 5486
rect 13832 5452 13836 5486
rect 13874 5452 13900 5486
rect 13900 5452 13908 5486
rect 13976 5452 13984 5486
rect 13984 5452 14010 5486
rect 14048 5452 14052 5486
rect 14052 5452 14082 5486
rect 14120 5452 14154 5486
rect 14192 5452 14222 5486
rect 14222 5452 14226 5486
rect 14264 5452 14290 5486
rect 14290 5452 14298 5486
rect 14366 5452 14374 5486
rect 14374 5452 14400 5486
rect 14438 5452 14442 5486
rect 14442 5452 14472 5486
rect 14510 5452 14544 5486
rect 14582 5452 14612 5486
rect 14612 5452 14616 5486
rect 14654 5452 14680 5486
rect 14680 5452 14688 5486
rect 14756 5452 14764 5486
rect 14764 5452 14790 5486
rect 14828 5452 14832 5486
rect 14832 5452 14862 5486
rect 14900 5452 14934 5486
rect 14972 5452 15002 5486
rect 15002 5452 15006 5486
rect 15044 5452 15070 5486
rect 15070 5452 15078 5486
rect 24614 5452 24648 5486
rect 24696 5452 24730 5486
rect 24788 5452 24796 5486
rect 24796 5452 24822 5486
rect 24860 5452 24864 5486
rect 24864 5452 24894 5486
rect 24932 5452 24966 5486
rect 25004 5452 25034 5486
rect 25034 5452 25038 5486
rect 25076 5452 25102 5486
rect 25102 5452 25110 5486
rect 25178 5452 25186 5486
rect 25186 5452 25212 5486
rect 25250 5452 25254 5486
rect 25254 5452 25284 5486
rect 25322 5452 25356 5486
rect 25394 5452 25424 5486
rect 25424 5452 25428 5486
rect 25466 5452 25492 5486
rect 25492 5452 25500 5486
rect 25568 5452 25576 5486
rect 25576 5452 25602 5486
rect 25640 5452 25644 5486
rect 25644 5452 25674 5486
rect 25712 5452 25746 5486
rect 25784 5452 25814 5486
rect 25814 5452 25818 5486
rect 25856 5452 25882 5486
rect 25882 5452 25890 5486
rect 25958 5452 25966 5486
rect 25966 5452 25992 5486
rect 26030 5452 26034 5486
rect 26034 5452 26064 5486
rect 26102 5452 26136 5486
rect 26174 5452 26204 5486
rect 26204 5452 26208 5486
rect 26246 5452 26272 5486
rect 26272 5452 26280 5486
rect 26348 5452 26356 5486
rect 26356 5452 26382 5486
rect 26420 5452 26424 5486
rect 26424 5452 26454 5486
rect 26492 5452 26526 5486
rect 26564 5452 26594 5486
rect 26594 5452 26598 5486
rect 26636 5452 26662 5486
rect 26662 5452 26670 5486
rect 13080 5319 13114 5353
rect 13210 5319 13244 5353
rect 13340 5319 13374 5353
rect 13470 5319 13504 5353
rect 13600 5319 13634 5353
rect 13730 5319 13764 5353
rect 13860 5319 13894 5353
rect 13990 5319 14024 5353
rect 14120 5319 14154 5353
rect 14250 5319 14284 5353
rect 14380 5319 14414 5353
rect 14510 5319 14544 5353
rect 14640 5319 14674 5353
rect 14770 5319 14804 5353
rect 14900 5319 14934 5353
rect 15030 5319 15064 5353
rect 24672 5319 24706 5353
rect 24802 5319 24836 5353
rect 24932 5319 24966 5353
rect 25062 5319 25096 5353
rect 25192 5319 25226 5353
rect 25322 5319 25356 5353
rect 25452 5319 25486 5353
rect 25582 5319 25616 5353
rect 25712 5319 25746 5353
rect 25842 5319 25876 5353
rect 25972 5319 26006 5353
rect 26102 5319 26136 5353
rect 26232 5319 26266 5353
rect 26362 5319 26396 5353
rect 26492 5319 26526 5353
rect 26622 5319 26656 5353
rect 13015 5190 13049 5224
rect 13015 5118 13049 5152
rect 13015 5046 13049 5080
rect 13015 4974 13049 5008
rect 13015 4902 13049 4936
rect 13145 5190 13179 5224
rect 13145 5118 13179 5152
rect 13145 5046 13179 5080
rect 13145 4974 13179 5008
rect 13145 4902 13179 4936
rect 13275 5190 13309 5224
rect 13275 5118 13309 5152
rect 13275 5046 13309 5080
rect 13275 4974 13309 5008
rect 13275 4902 13309 4936
rect 13405 5190 13439 5224
rect 13405 5118 13439 5152
rect 13405 5046 13439 5080
rect 13405 4974 13439 5008
rect 13405 4902 13439 4936
rect 13535 5190 13569 5224
rect 13535 5118 13569 5152
rect 13535 5046 13569 5080
rect 13535 4974 13569 5008
rect 13535 4902 13569 4936
rect 13665 5190 13699 5224
rect 13665 5118 13699 5152
rect 13665 5046 13699 5080
rect 13665 4974 13699 5008
rect 13665 4902 13699 4936
rect 13795 5190 13829 5224
rect 13795 5118 13829 5152
rect 13795 5046 13829 5080
rect 13795 4974 13829 5008
rect 13795 4902 13829 4936
rect 13925 5190 13959 5224
rect 13925 5118 13959 5152
rect 13925 5046 13959 5080
rect 13925 4974 13959 5008
rect 13925 4902 13959 4936
rect 14055 5190 14089 5224
rect 14055 5118 14089 5152
rect 14055 5046 14089 5080
rect 14055 4974 14089 5008
rect 14055 4902 14089 4936
rect 14185 5190 14219 5224
rect 14185 5118 14219 5152
rect 14185 5046 14219 5080
rect 14185 4974 14219 5008
rect 14185 4902 14219 4936
rect 14315 5190 14349 5224
rect 14315 5118 14349 5152
rect 14315 5046 14349 5080
rect 14315 4974 14349 5008
rect 14315 4902 14349 4936
rect 14445 5190 14479 5224
rect 14445 5118 14479 5152
rect 14445 5046 14479 5080
rect 14445 4974 14479 5008
rect 14445 4902 14479 4936
rect 14575 5190 14609 5224
rect 14575 5118 14609 5152
rect 14575 5046 14609 5080
rect 14575 4974 14609 5008
rect 14575 4902 14609 4936
rect 14705 5190 14739 5224
rect 14705 5118 14739 5152
rect 14705 5046 14739 5080
rect 14705 4974 14739 5008
rect 14705 4902 14739 4936
rect 14835 5190 14869 5224
rect 14835 5118 14869 5152
rect 14835 5046 14869 5080
rect 14835 4974 14869 5008
rect 14835 4902 14869 4936
rect 14965 5190 14999 5224
rect 14965 5118 14999 5152
rect 14965 5046 14999 5080
rect 14965 4974 14999 5008
rect 14965 4902 14999 4936
rect 15095 5190 15129 5224
rect 15095 5118 15129 5152
rect 15095 5046 15129 5080
rect 15095 4974 15129 5008
rect 15095 4902 15129 4936
rect 24607 5190 24641 5224
rect 24607 5118 24641 5152
rect 24607 5046 24641 5080
rect 24607 4974 24641 5008
rect 15315 4881 15319 4915
rect 15319 4881 15349 4915
rect 15387 4881 15421 4915
rect 15459 4881 15489 4915
rect 15489 4881 15493 4915
rect 24607 4902 24641 4936
rect 24737 5190 24771 5224
rect 24737 5118 24771 5152
rect 24737 5046 24771 5080
rect 24737 4974 24771 5008
rect 24737 4902 24771 4936
rect 24867 5190 24901 5224
rect 24867 5118 24901 5152
rect 24867 5046 24901 5080
rect 24867 4974 24901 5008
rect 24867 4902 24901 4936
rect 24997 5190 25031 5224
rect 24997 5118 25031 5152
rect 24997 5046 25031 5080
rect 24997 4974 25031 5008
rect 24997 4902 25031 4936
rect 25127 5190 25161 5224
rect 25127 5118 25161 5152
rect 25127 5046 25161 5080
rect 25127 4974 25161 5008
rect 25127 4902 25161 4936
rect 25257 5190 25291 5224
rect 25257 5118 25291 5152
rect 25257 5046 25291 5080
rect 25257 4974 25291 5008
rect 25257 4902 25291 4936
rect 25387 5190 25421 5224
rect 25387 5118 25421 5152
rect 25387 5046 25421 5080
rect 25387 4974 25421 5008
rect 25387 4902 25421 4936
rect 25517 5190 25551 5224
rect 25517 5118 25551 5152
rect 25517 5046 25551 5080
rect 25517 4974 25551 5008
rect 25517 4902 25551 4936
rect 25647 5190 25681 5224
rect 25647 5118 25681 5152
rect 25647 5046 25681 5080
rect 25647 4974 25681 5008
rect 25647 4902 25681 4936
rect 25777 5190 25811 5224
rect 25777 5118 25811 5152
rect 25777 5046 25811 5080
rect 25777 4974 25811 5008
rect 25777 4902 25811 4936
rect 25907 5190 25941 5224
rect 25907 5118 25941 5152
rect 25907 5046 25941 5080
rect 25907 4974 25941 5008
rect 25907 4902 25941 4936
rect 26037 5190 26071 5224
rect 26037 5118 26071 5152
rect 26037 5046 26071 5080
rect 26037 4974 26071 5008
rect 26037 4902 26071 4936
rect 26167 5190 26201 5224
rect 26167 5118 26201 5152
rect 26167 5046 26201 5080
rect 26167 4974 26201 5008
rect 26167 4902 26201 4936
rect 26297 5190 26331 5224
rect 26297 5118 26331 5152
rect 26297 5046 26331 5080
rect 26297 4974 26331 5008
rect 26297 4902 26331 4936
rect 26427 5190 26461 5224
rect 26427 5118 26461 5152
rect 26427 5046 26461 5080
rect 26427 4974 26461 5008
rect 26427 4902 26461 4936
rect 26557 5190 26591 5224
rect 26557 5118 26591 5152
rect 26557 5046 26591 5080
rect 26557 4974 26591 5008
rect 26557 4902 26591 4936
rect 26687 5190 26721 5224
rect 26687 5118 26721 5152
rect 26687 5046 26721 5080
rect 26687 4974 26721 5008
rect 26687 4902 26721 4936
rect 26907 4881 26911 4915
rect 26911 4881 26941 4915
rect 26979 4881 27013 4915
rect 27051 4881 27081 4915
rect 27081 4881 27085 4915
rect 15402 4790 15404 4824
rect 15404 4790 15436 4824
rect 15474 4790 15506 4824
rect 15506 4790 15508 4824
rect 26994 4790 26996 4824
rect 26996 4790 27028 4824
rect 27066 4790 27098 4824
rect 27098 4790 27100 4824
rect 13275 4642 13309 4676
rect 13275 4570 13309 4604
rect 13275 4498 13309 4532
rect 13275 4426 13309 4460
rect 13275 4354 13309 4388
rect 13405 4642 13439 4676
rect 13405 4570 13439 4604
rect 13405 4498 13439 4532
rect 13405 4426 13439 4460
rect 13405 4354 13439 4388
rect 13665 4642 13699 4676
rect 13665 4570 13699 4604
rect 13665 4498 13699 4532
rect 13665 4426 13699 4460
rect 13665 4354 13699 4388
rect 13795 4642 13829 4676
rect 13795 4570 13829 4604
rect 13795 4498 13829 4532
rect 13795 4426 13829 4460
rect 13795 4354 13829 4388
rect 14055 4642 14089 4676
rect 14055 4570 14089 4604
rect 14055 4498 14089 4532
rect 14055 4426 14089 4460
rect 14055 4354 14089 4388
rect 14185 4642 14219 4676
rect 14185 4570 14219 4604
rect 14185 4498 14219 4532
rect 14185 4426 14219 4460
rect 14185 4354 14219 4388
rect 14445 4642 14479 4676
rect 14445 4570 14479 4604
rect 14445 4498 14479 4532
rect 14445 4426 14479 4460
rect 14445 4354 14479 4388
rect 14575 4642 14609 4676
rect 14575 4570 14609 4604
rect 14575 4498 14609 4532
rect 14575 4426 14609 4460
rect 14575 4354 14609 4388
rect 14835 4642 14869 4676
rect 14835 4570 14869 4604
rect 14835 4498 14869 4532
rect 14835 4426 14869 4460
rect 14835 4354 14869 4388
rect 14965 4642 14999 4676
rect 14965 4570 14999 4604
rect 14965 4498 14999 4532
rect 14965 4426 14999 4460
rect 14965 4354 14999 4388
rect 15209 4642 15243 4676
rect 15209 4570 15243 4604
rect 15209 4498 15243 4532
rect 15209 4426 15243 4460
rect 15209 4354 15243 4388
rect 15299 4642 15333 4676
rect 15299 4570 15333 4604
rect 15299 4498 15333 4532
rect 15299 4426 15333 4460
rect 15299 4354 15333 4388
rect 15389 4642 15423 4676
rect 15389 4570 15423 4604
rect 15389 4498 15423 4532
rect 15389 4426 15423 4460
rect 15389 4354 15423 4388
rect 15479 4642 15513 4676
rect 15479 4570 15513 4604
rect 15479 4498 15513 4532
rect 15479 4426 15513 4460
rect 15479 4354 15513 4388
rect 15569 4642 15603 4676
rect 15569 4570 15603 4604
rect 15569 4498 15603 4532
rect 15569 4426 15603 4460
rect 15569 4354 15603 4388
rect 24867 4642 24901 4676
rect 24867 4570 24901 4604
rect 24867 4498 24901 4532
rect 24867 4426 24901 4460
rect 24867 4354 24901 4388
rect 24997 4642 25031 4676
rect 24997 4570 25031 4604
rect 24997 4498 25031 4532
rect 24997 4426 25031 4460
rect 24997 4354 25031 4388
rect 25257 4642 25291 4676
rect 25257 4570 25291 4604
rect 25257 4498 25291 4532
rect 25257 4426 25291 4460
rect 25257 4354 25291 4388
rect 25387 4642 25421 4676
rect 25387 4570 25421 4604
rect 25387 4498 25421 4532
rect 25387 4426 25421 4460
rect 25387 4354 25421 4388
rect 25647 4642 25681 4676
rect 25647 4570 25681 4604
rect 25647 4498 25681 4532
rect 25647 4426 25681 4460
rect 25647 4354 25681 4388
rect 25777 4642 25811 4676
rect 25777 4570 25811 4604
rect 25777 4498 25811 4532
rect 25777 4426 25811 4460
rect 25777 4354 25811 4388
rect 26037 4642 26071 4676
rect 26037 4570 26071 4604
rect 26037 4498 26071 4532
rect 26037 4426 26071 4460
rect 26037 4354 26071 4388
rect 26167 4642 26201 4676
rect 26167 4570 26201 4604
rect 26167 4498 26201 4532
rect 26167 4426 26201 4460
rect 26167 4354 26201 4388
rect 26427 4642 26461 4676
rect 26427 4570 26461 4604
rect 26427 4498 26461 4532
rect 26427 4426 26461 4460
rect 26427 4354 26461 4388
rect 26557 4642 26591 4676
rect 26557 4570 26591 4604
rect 26557 4498 26591 4532
rect 26557 4426 26591 4460
rect 26557 4354 26591 4388
rect 26801 4642 26835 4676
rect 26801 4570 26835 4604
rect 26801 4498 26835 4532
rect 26801 4426 26835 4460
rect 26801 4354 26835 4388
rect 26891 4642 26925 4676
rect 26891 4570 26925 4604
rect 26891 4498 26925 4532
rect 26891 4426 26925 4460
rect 26891 4354 26925 4388
rect 26981 4642 27015 4676
rect 26981 4570 27015 4604
rect 26981 4498 27015 4532
rect 26981 4426 27015 4460
rect 26981 4354 27015 4388
rect 27071 4642 27105 4676
rect 27071 4570 27105 4604
rect 27071 4498 27105 4532
rect 27071 4426 27105 4460
rect 27071 4354 27105 4388
rect 27161 4642 27195 4676
rect 27161 4570 27195 4604
rect 27161 4498 27195 4532
rect 27161 4426 27195 4460
rect 27161 4354 27195 4388
rect 13244 4074 13278 4108
rect 13634 4074 13668 4108
rect 14024 4074 14058 4108
rect 14414 4074 14448 4108
rect 14804 4074 14838 4108
rect 15249 4074 15283 4108
rect 24836 4074 24870 4108
rect 25226 4074 25260 4108
rect 25616 4074 25650 4108
rect 26006 4074 26040 4108
rect 26396 4074 26430 4108
rect 26841 4074 26875 4108
rect 13860 3917 13894 3951
rect 14640 3917 14674 3951
rect 25452 3917 25486 3951
rect 26232 3917 26266 3951
rect 13275 3786 13309 3820
rect 13275 3714 13309 3748
rect 13405 3786 13439 3820
rect 13405 3714 13439 3748
rect 13535 3786 13569 3820
rect 13535 3714 13569 3748
rect 13665 3786 13699 3820
rect 13665 3714 13699 3748
rect 13795 3786 13829 3820
rect 13795 3714 13829 3748
rect 13925 3786 13959 3820
rect 13925 3714 13959 3748
rect 14055 3786 14089 3820
rect 14055 3714 14089 3748
rect 14185 3786 14219 3820
rect 14185 3714 14219 3748
rect 14315 3786 14349 3820
rect 14315 3714 14349 3748
rect 14445 3786 14479 3820
rect 14445 3714 14479 3748
rect 14575 3786 14609 3820
rect 14575 3714 14609 3748
rect 14705 3786 14739 3820
rect 14705 3714 14739 3748
rect 14835 3786 14869 3820
rect 14835 3714 14869 3748
rect 14965 3786 14999 3820
rect 14965 3714 14999 3748
rect 15095 3786 15129 3820
rect 15095 3714 15129 3748
rect 15209 3786 15243 3820
rect 15209 3714 15243 3748
rect 15299 3786 15333 3820
rect 15299 3714 15333 3748
rect 15389 3786 15423 3820
rect 15389 3714 15423 3748
rect 15479 3786 15513 3820
rect 15479 3714 15513 3748
rect 15569 3786 15603 3820
rect 15569 3714 15603 3748
rect 24867 3786 24901 3820
rect 24867 3714 24901 3748
rect 24997 3786 25031 3820
rect 24997 3714 25031 3748
rect 25127 3786 25161 3820
rect 25127 3714 25161 3748
rect 25257 3786 25291 3820
rect 25257 3714 25291 3748
rect 25387 3786 25421 3820
rect 25387 3714 25421 3748
rect 25517 3786 25551 3820
rect 25517 3714 25551 3748
rect 25647 3786 25681 3820
rect 25647 3714 25681 3748
rect 25777 3786 25811 3820
rect 25777 3714 25811 3748
rect 25907 3786 25941 3820
rect 25907 3714 25941 3748
rect 26037 3786 26071 3820
rect 26037 3714 26071 3748
rect 26167 3786 26201 3820
rect 26167 3714 26201 3748
rect 26297 3786 26331 3820
rect 26297 3714 26331 3748
rect 26427 3786 26461 3820
rect 26427 3714 26461 3748
rect 26557 3786 26591 3820
rect 26557 3714 26591 3748
rect 26687 3786 26721 3820
rect 26687 3714 26721 3748
rect 26801 3786 26835 3820
rect 26801 3714 26835 3748
rect 26891 3786 26925 3820
rect 26891 3714 26925 3748
rect 26981 3786 27015 3820
rect 26981 3714 27015 3748
rect 27071 3786 27105 3820
rect 27071 3714 27105 3748
rect 27161 3786 27195 3820
rect 27161 3714 27195 3748
rect 15318 3545 15322 3579
rect 15322 3545 15352 3579
rect 15390 3545 15424 3579
rect 15462 3545 15492 3579
rect 15492 3545 15496 3579
rect 26910 3545 26914 3579
rect 26914 3545 26944 3579
rect 26982 3545 27016 3579
rect 27054 3545 27084 3579
rect 27084 3545 27088 3579
rect 13015 3438 13049 3472
rect 13015 3366 13049 3400
rect 13145 3438 13179 3472
rect 13145 3366 13179 3400
rect 13275 3438 13309 3472
rect 13275 3366 13309 3400
rect 13405 3438 13439 3472
rect 13405 3366 13439 3400
rect 13535 3438 13569 3472
rect 13535 3366 13569 3400
rect 13665 3438 13699 3472
rect 13665 3366 13699 3400
rect 13795 3438 13829 3472
rect 13795 3366 13829 3400
rect 13925 3438 13959 3472
rect 13925 3366 13959 3400
rect 14055 3438 14089 3472
rect 14055 3366 14089 3400
rect 14185 3438 14219 3472
rect 14185 3366 14219 3400
rect 14315 3438 14349 3472
rect 14315 3366 14349 3400
rect 14445 3438 14479 3472
rect 14445 3366 14479 3400
rect 14575 3438 14609 3472
rect 14575 3366 14609 3400
rect 14705 3438 14739 3472
rect 14705 3366 14739 3400
rect 14835 3438 14869 3472
rect 14835 3366 14869 3400
rect 14965 3438 14999 3472
rect 14965 3366 14999 3400
rect 15095 3438 15129 3472
rect 15095 3366 15129 3400
rect 24607 3438 24641 3472
rect 24607 3366 24641 3400
rect 24737 3438 24771 3472
rect 24737 3366 24771 3400
rect 24867 3438 24901 3472
rect 24867 3366 24901 3400
rect 24997 3438 25031 3472
rect 24997 3366 25031 3400
rect 25127 3438 25161 3472
rect 25127 3366 25161 3400
rect 25257 3438 25291 3472
rect 25257 3366 25291 3400
rect 25387 3438 25421 3472
rect 25387 3366 25421 3400
rect 25517 3438 25551 3472
rect 25517 3366 25551 3400
rect 25647 3438 25681 3472
rect 25647 3366 25681 3400
rect 25777 3438 25811 3472
rect 25777 3366 25811 3400
rect 25907 3438 25941 3472
rect 25907 3366 25941 3400
rect 26037 3438 26071 3472
rect 26037 3366 26071 3400
rect 26167 3438 26201 3472
rect 26167 3366 26201 3400
rect 26297 3438 26331 3472
rect 26297 3366 26331 3400
rect 26427 3438 26461 3472
rect 26427 3366 26461 3400
rect 26557 3438 26591 3472
rect 26557 3366 26591 3400
rect 26687 3438 26721 3472
rect 26687 3366 26721 3400
rect 13012 3229 13046 3263
rect 13210 3229 13244 3263
rect 13340 3229 13374 3263
rect 13470 3229 13504 3263
rect 13600 3229 13634 3263
rect 13730 3229 13764 3263
rect 13860 3229 13894 3263
rect 13990 3229 14024 3263
rect 14120 3229 14154 3263
rect 14250 3229 14284 3263
rect 14380 3229 14414 3263
rect 14510 3229 14544 3263
rect 14640 3229 14674 3263
rect 14770 3229 14804 3263
rect 14900 3229 14934 3263
rect 15030 3229 15064 3263
rect 24604 3229 24638 3263
rect 24802 3229 24836 3263
rect 24932 3229 24966 3263
rect 25062 3229 25096 3263
rect 25192 3229 25226 3263
rect 25322 3229 25356 3263
rect 25452 3229 25486 3263
rect 25582 3229 25616 3263
rect 25712 3229 25746 3263
rect 25842 3229 25876 3263
rect 25972 3229 26006 3263
rect 26102 3229 26136 3263
rect 26232 3229 26266 3263
rect 26362 3229 26396 3263
rect 26492 3229 26526 3263
rect 26622 3229 26656 3263
rect 13022 3096 13056 3130
rect 13104 3096 13138 3130
rect 13196 3096 13204 3130
rect 13204 3096 13230 3130
rect 13268 3096 13272 3130
rect 13272 3096 13302 3130
rect 13340 3096 13374 3130
rect 13412 3096 13442 3130
rect 13442 3096 13446 3130
rect 13484 3096 13510 3130
rect 13510 3096 13518 3130
rect 13586 3096 13594 3130
rect 13594 3096 13620 3130
rect 13658 3096 13662 3130
rect 13662 3096 13692 3130
rect 13730 3096 13764 3130
rect 13802 3096 13832 3130
rect 13832 3096 13836 3130
rect 13874 3096 13900 3130
rect 13900 3096 13908 3130
rect 13976 3096 13984 3130
rect 13984 3096 14010 3130
rect 14048 3096 14052 3130
rect 14052 3096 14082 3130
rect 14120 3096 14154 3130
rect 14192 3096 14222 3130
rect 14222 3096 14226 3130
rect 14264 3096 14290 3130
rect 14290 3096 14298 3130
rect 14366 3096 14374 3130
rect 14374 3096 14400 3130
rect 14438 3096 14442 3130
rect 14442 3096 14472 3130
rect 14510 3096 14544 3130
rect 14582 3096 14612 3130
rect 14612 3096 14616 3130
rect 14654 3096 14680 3130
rect 14680 3096 14688 3130
rect 14756 3096 14764 3130
rect 14764 3096 14790 3130
rect 14828 3096 14832 3130
rect 14832 3096 14862 3130
rect 14900 3096 14934 3130
rect 14972 3096 15002 3130
rect 15002 3096 15006 3130
rect 15044 3096 15070 3130
rect 15070 3096 15078 3130
rect 15146 3096 15154 3130
rect 15154 3096 15180 3130
rect 15218 3096 15222 3130
rect 15222 3096 15252 3130
rect 15290 3096 15324 3130
rect 15362 3096 15392 3130
rect 15392 3096 15396 3130
rect 15434 3096 15460 3130
rect 15460 3096 15468 3130
rect 24614 3096 24648 3130
rect 24696 3096 24730 3130
rect 24788 3096 24796 3130
rect 24796 3096 24822 3130
rect 24860 3096 24864 3130
rect 24864 3096 24894 3130
rect 24932 3096 24966 3130
rect 25004 3096 25034 3130
rect 25034 3096 25038 3130
rect 25076 3096 25102 3130
rect 25102 3096 25110 3130
rect 25178 3096 25186 3130
rect 25186 3096 25212 3130
rect 25250 3096 25254 3130
rect 25254 3096 25284 3130
rect 25322 3096 25356 3130
rect 25394 3096 25424 3130
rect 25424 3096 25428 3130
rect 25466 3096 25492 3130
rect 25492 3096 25500 3130
rect 25568 3096 25576 3130
rect 25576 3096 25602 3130
rect 25640 3096 25644 3130
rect 25644 3096 25674 3130
rect 25712 3096 25746 3130
rect 25784 3096 25814 3130
rect 25814 3096 25818 3130
rect 25856 3096 25882 3130
rect 25882 3096 25890 3130
rect 25958 3096 25966 3130
rect 25966 3096 25992 3130
rect 26030 3096 26034 3130
rect 26034 3096 26064 3130
rect 26102 3096 26136 3130
rect 26174 3096 26204 3130
rect 26204 3096 26208 3130
rect 26246 3096 26272 3130
rect 26272 3096 26280 3130
rect 26348 3096 26356 3130
rect 26356 3096 26382 3130
rect 26420 3096 26424 3130
rect 26424 3096 26454 3130
rect 26492 3096 26526 3130
rect 26564 3096 26594 3130
rect 26594 3096 26598 3130
rect 26636 3096 26662 3130
rect 26662 3096 26670 3130
rect 26738 3096 26746 3130
rect 26746 3096 26772 3130
rect 26810 3096 26814 3130
rect 26814 3096 26844 3130
rect 26882 3096 26916 3130
rect 26954 3096 26984 3130
rect 26984 3096 26988 3130
rect 27026 3096 27052 3130
rect 27052 3096 27060 3130
rect 13210 2963 13244 2997
rect 13340 2963 13374 2997
rect 13470 2963 13504 2997
rect 13600 2963 13634 2997
rect 13730 2963 13764 2997
rect 13860 2963 13894 2997
rect 13990 2963 14024 2997
rect 14120 2963 14154 2997
rect 14250 2963 14284 2997
rect 14380 2963 14414 2997
rect 14510 2963 14544 2997
rect 14640 2963 14674 2997
rect 14770 2963 14804 2997
rect 14900 2963 14934 2997
rect 15030 2963 15064 2997
rect 15160 2963 15194 2997
rect 15290 2963 15324 2997
rect 15420 2963 15454 2997
rect 24802 2963 24836 2997
rect 24932 2963 24966 2997
rect 25062 2963 25096 2997
rect 25192 2963 25226 2997
rect 25322 2963 25356 2997
rect 25452 2963 25486 2997
rect 25582 2963 25616 2997
rect 25712 2963 25746 2997
rect 25842 2963 25876 2997
rect 25972 2963 26006 2997
rect 26102 2963 26136 2997
rect 26232 2963 26266 2997
rect 26362 2963 26396 2997
rect 26492 2963 26526 2997
rect 26622 2963 26656 2997
rect 26752 2963 26786 2997
rect 26882 2963 26916 2997
rect 27012 2963 27046 2997
rect 13145 2826 13179 2860
rect 13145 2754 13179 2788
rect 13275 2826 13309 2860
rect 13275 2754 13309 2788
rect 13405 2826 13439 2860
rect 13405 2754 13439 2788
rect 13535 2826 13569 2860
rect 13535 2754 13569 2788
rect 13665 2826 13699 2860
rect 13665 2754 13699 2788
rect 13795 2826 13829 2860
rect 13795 2754 13829 2788
rect 13925 2826 13959 2860
rect 13925 2754 13959 2788
rect 14055 2826 14089 2860
rect 14055 2754 14089 2788
rect 14185 2826 14219 2860
rect 14185 2754 14219 2788
rect 14315 2826 14349 2860
rect 14315 2754 14349 2788
rect 14445 2826 14479 2860
rect 14445 2754 14479 2788
rect 14575 2826 14609 2860
rect 14575 2754 14609 2788
rect 14705 2826 14739 2860
rect 14705 2754 14739 2788
rect 14835 2826 14869 2860
rect 14835 2754 14869 2788
rect 14965 2826 14999 2860
rect 14965 2754 14999 2788
rect 15095 2826 15129 2860
rect 15095 2754 15129 2788
rect 15225 2826 15259 2860
rect 15225 2754 15259 2788
rect 15355 2826 15389 2860
rect 15355 2754 15389 2788
rect 15485 2826 15519 2860
rect 15485 2754 15519 2788
rect 24737 2826 24771 2860
rect 24737 2754 24771 2788
rect 24867 2826 24901 2860
rect 24867 2754 24901 2788
rect 24997 2826 25031 2860
rect 24997 2754 25031 2788
rect 25127 2826 25161 2860
rect 25127 2754 25161 2788
rect 25257 2826 25291 2860
rect 25257 2754 25291 2788
rect 25387 2826 25421 2860
rect 25387 2754 25421 2788
rect 25517 2826 25551 2860
rect 25517 2754 25551 2788
rect 25647 2826 25681 2860
rect 25647 2754 25681 2788
rect 25777 2826 25811 2860
rect 25777 2754 25811 2788
rect 25907 2826 25941 2860
rect 25907 2754 25941 2788
rect 26037 2826 26071 2860
rect 26037 2754 26071 2788
rect 26167 2826 26201 2860
rect 26167 2754 26201 2788
rect 26297 2826 26331 2860
rect 26297 2754 26331 2788
rect 26427 2826 26461 2860
rect 26427 2754 26461 2788
rect 26557 2826 26591 2860
rect 26557 2754 26591 2788
rect 26687 2826 26721 2860
rect 26687 2754 26721 2788
rect 26817 2826 26851 2860
rect 26817 2754 26851 2788
rect 26947 2826 26981 2860
rect 26947 2754 26981 2788
rect 27077 2826 27111 2860
rect 27077 2754 27111 2788
rect 13145 2478 13179 2512
rect 13145 2406 13179 2440
rect 13275 2478 13309 2512
rect 13275 2406 13309 2440
rect 13405 2478 13439 2512
rect 13405 2406 13439 2440
rect 13535 2478 13569 2512
rect 13535 2406 13569 2440
rect 13665 2478 13699 2512
rect 13665 2406 13699 2440
rect 13795 2478 13829 2512
rect 13795 2406 13829 2440
rect 13925 2478 13959 2512
rect 13925 2406 13959 2440
rect 14055 2478 14089 2512
rect 14055 2406 14089 2440
rect 14185 2478 14219 2512
rect 14185 2406 14219 2440
rect 14315 2478 14349 2512
rect 14315 2406 14349 2440
rect 14445 2478 14479 2512
rect 14445 2406 14479 2440
rect 14575 2478 14609 2512
rect 14575 2406 14609 2440
rect 14705 2478 14739 2512
rect 14705 2406 14739 2440
rect 14835 2478 14869 2512
rect 14835 2406 14869 2440
rect 14965 2478 14999 2512
rect 14965 2406 14999 2440
rect 15095 2478 15129 2512
rect 15095 2406 15129 2440
rect 15225 2478 15259 2512
rect 15225 2406 15259 2440
rect 15355 2478 15389 2512
rect 15355 2406 15389 2440
rect 24737 2478 24771 2512
rect 24737 2406 24771 2440
rect 24867 2478 24901 2512
rect 24867 2406 24901 2440
rect 24997 2478 25031 2512
rect 24997 2406 25031 2440
rect 25127 2478 25161 2512
rect 25127 2406 25161 2440
rect 25257 2478 25291 2512
rect 25257 2406 25291 2440
rect 25387 2478 25421 2512
rect 25387 2406 25421 2440
rect 25517 2478 25551 2512
rect 25517 2406 25551 2440
rect 25647 2478 25681 2512
rect 25647 2406 25681 2440
rect 25777 2478 25811 2512
rect 25777 2406 25811 2440
rect 25907 2478 25941 2512
rect 25907 2406 25941 2440
rect 26037 2478 26071 2512
rect 26037 2406 26071 2440
rect 26167 2478 26201 2512
rect 26167 2406 26201 2440
rect 26297 2478 26331 2512
rect 26297 2406 26331 2440
rect 26427 2478 26461 2512
rect 26427 2406 26461 2440
rect 26557 2478 26591 2512
rect 26557 2406 26591 2440
rect 26687 2478 26721 2512
rect 26687 2406 26721 2440
rect 26817 2478 26851 2512
rect 26817 2406 26851 2440
rect 26947 2478 26981 2512
rect 26947 2406 26981 2440
rect 13210 2275 13244 2309
rect 13600 2275 13634 2309
rect 14380 2275 14414 2309
rect 15160 2275 15194 2309
rect 24802 2275 24836 2309
rect 25192 2275 25226 2309
rect 25972 2275 26006 2309
rect 26752 2275 26786 2309
rect 13436 2118 13470 2152
rect 13826 2118 13860 2152
rect 14216 2118 14250 2152
rect 14606 2118 14640 2152
rect 14996 2118 15030 2152
rect 15386 2118 15420 2152
rect 25028 2118 25062 2152
rect 25418 2118 25452 2152
rect 25808 2118 25842 2152
rect 26198 2118 26232 2152
rect 26588 2118 26622 2152
rect 26978 2118 27012 2152
rect 13275 1838 13309 1872
rect 13275 1766 13309 1800
rect 13275 1694 13309 1728
rect 13275 1622 13309 1656
rect 13275 1550 13309 1584
rect 13405 1838 13439 1872
rect 13405 1766 13439 1800
rect 13405 1694 13439 1728
rect 13405 1622 13439 1656
rect 13405 1550 13439 1584
rect 13665 1838 13699 1872
rect 13665 1766 13699 1800
rect 13665 1694 13699 1728
rect 13665 1622 13699 1656
rect 13665 1550 13699 1584
rect 13795 1838 13829 1872
rect 13795 1766 13829 1800
rect 13795 1694 13829 1728
rect 13795 1622 13829 1656
rect 13795 1550 13829 1584
rect 14055 1838 14089 1872
rect 14055 1766 14089 1800
rect 14055 1694 14089 1728
rect 14055 1622 14089 1656
rect 14055 1550 14089 1584
rect 14185 1838 14219 1872
rect 14185 1766 14219 1800
rect 14185 1694 14219 1728
rect 14185 1622 14219 1656
rect 14185 1550 14219 1584
rect 14445 1838 14479 1872
rect 14445 1766 14479 1800
rect 14445 1694 14479 1728
rect 14445 1622 14479 1656
rect 14445 1550 14479 1584
rect 14575 1838 14609 1872
rect 14575 1766 14609 1800
rect 14575 1694 14609 1728
rect 14575 1622 14609 1656
rect 14575 1550 14609 1584
rect 14835 1838 14869 1872
rect 14835 1766 14869 1800
rect 14835 1694 14869 1728
rect 14835 1622 14869 1656
rect 14835 1550 14869 1584
rect 14965 1838 14999 1872
rect 14965 1766 14999 1800
rect 14965 1694 14999 1728
rect 14965 1622 14999 1656
rect 14965 1550 14999 1584
rect 15225 1838 15259 1872
rect 15225 1766 15259 1800
rect 15225 1694 15259 1728
rect 15225 1622 15259 1656
rect 15225 1550 15259 1584
rect 15355 1838 15389 1872
rect 15355 1766 15389 1800
rect 15355 1694 15389 1728
rect 15355 1622 15389 1656
rect 15355 1550 15389 1584
rect 24867 1838 24901 1872
rect 24867 1766 24901 1800
rect 24867 1694 24901 1728
rect 24867 1622 24901 1656
rect 24867 1550 24901 1584
rect 24997 1838 25031 1872
rect 24997 1766 25031 1800
rect 24997 1694 25031 1728
rect 24997 1622 25031 1656
rect 24997 1550 25031 1584
rect 25257 1838 25291 1872
rect 25257 1766 25291 1800
rect 25257 1694 25291 1728
rect 25257 1622 25291 1656
rect 25257 1550 25291 1584
rect 25387 1838 25421 1872
rect 25387 1766 25421 1800
rect 25387 1694 25421 1728
rect 25387 1622 25421 1656
rect 25387 1550 25421 1584
rect 25647 1838 25681 1872
rect 25647 1766 25681 1800
rect 25647 1694 25681 1728
rect 25647 1622 25681 1656
rect 25647 1550 25681 1584
rect 25777 1838 25811 1872
rect 25777 1766 25811 1800
rect 25777 1694 25811 1728
rect 25777 1622 25811 1656
rect 25777 1550 25811 1584
rect 26037 1838 26071 1872
rect 26037 1766 26071 1800
rect 26037 1694 26071 1728
rect 26037 1622 26071 1656
rect 26037 1550 26071 1584
rect 26167 1838 26201 1872
rect 26167 1766 26201 1800
rect 26167 1694 26201 1728
rect 26167 1622 26201 1656
rect 26167 1550 26201 1584
rect 26427 1838 26461 1872
rect 26427 1766 26461 1800
rect 26427 1694 26461 1728
rect 26427 1622 26461 1656
rect 26427 1550 26461 1584
rect 26557 1838 26591 1872
rect 26557 1766 26591 1800
rect 26557 1694 26591 1728
rect 26557 1622 26591 1656
rect 26557 1550 26591 1584
rect 26817 1838 26851 1872
rect 26817 1766 26851 1800
rect 26817 1694 26851 1728
rect 26817 1622 26851 1656
rect 26817 1550 26851 1584
rect 26947 1838 26981 1872
rect 26947 1766 26981 1800
rect 26947 1694 26981 1728
rect 26947 1622 26981 1656
rect 26947 1550 26981 1584
rect 13145 1290 13179 1324
rect 13145 1218 13179 1252
rect 13145 1146 13179 1180
rect 13145 1074 13179 1108
rect 13145 1002 13179 1036
rect 13275 1290 13309 1324
rect 13275 1218 13309 1252
rect 13275 1146 13309 1180
rect 13275 1074 13309 1108
rect 13275 1002 13309 1036
rect 13405 1290 13439 1324
rect 13405 1218 13439 1252
rect 13405 1146 13439 1180
rect 13405 1074 13439 1108
rect 13405 1002 13439 1036
rect 13535 1290 13569 1324
rect 13535 1218 13569 1252
rect 13535 1146 13569 1180
rect 13535 1074 13569 1108
rect 13535 1002 13569 1036
rect 13665 1290 13699 1324
rect 13665 1218 13699 1252
rect 13665 1146 13699 1180
rect 13665 1074 13699 1108
rect 13665 1002 13699 1036
rect 13795 1290 13829 1324
rect 13795 1218 13829 1252
rect 13795 1146 13829 1180
rect 13795 1074 13829 1108
rect 13795 1002 13829 1036
rect 13925 1290 13959 1324
rect 13925 1218 13959 1252
rect 13925 1146 13959 1180
rect 13925 1074 13959 1108
rect 13925 1002 13959 1036
rect 14055 1290 14089 1324
rect 14055 1218 14089 1252
rect 14055 1146 14089 1180
rect 14055 1074 14089 1108
rect 14055 1002 14089 1036
rect 14185 1290 14219 1324
rect 14185 1218 14219 1252
rect 14185 1146 14219 1180
rect 14185 1074 14219 1108
rect 14185 1002 14219 1036
rect 14315 1290 14349 1324
rect 14315 1218 14349 1252
rect 14315 1146 14349 1180
rect 14315 1074 14349 1108
rect 14315 1002 14349 1036
rect 14445 1290 14479 1324
rect 14445 1218 14479 1252
rect 14445 1146 14479 1180
rect 14445 1074 14479 1108
rect 14445 1002 14479 1036
rect 14575 1290 14609 1324
rect 14575 1218 14609 1252
rect 14575 1146 14609 1180
rect 14575 1074 14609 1108
rect 14575 1002 14609 1036
rect 14705 1290 14739 1324
rect 14705 1218 14739 1252
rect 14705 1146 14739 1180
rect 14705 1074 14739 1108
rect 14705 1002 14739 1036
rect 14835 1290 14869 1324
rect 14835 1218 14869 1252
rect 14835 1146 14869 1180
rect 14835 1074 14869 1108
rect 14835 1002 14869 1036
rect 14965 1290 14999 1324
rect 14965 1218 14999 1252
rect 14965 1146 14999 1180
rect 14965 1074 14999 1108
rect 14965 1002 14999 1036
rect 15095 1290 15129 1324
rect 15095 1218 15129 1252
rect 15095 1146 15129 1180
rect 15095 1074 15129 1108
rect 15095 1002 15129 1036
rect 15225 1290 15259 1324
rect 15225 1218 15259 1252
rect 15225 1146 15259 1180
rect 15225 1074 15259 1108
rect 15225 1002 15259 1036
rect 15355 1290 15389 1324
rect 15355 1218 15389 1252
rect 15355 1146 15389 1180
rect 15355 1074 15389 1108
rect 15355 1002 15389 1036
rect 15485 1290 15519 1324
rect 15485 1218 15519 1252
rect 15485 1146 15519 1180
rect 15485 1074 15519 1108
rect 15485 1002 15519 1036
rect 24737 1290 24771 1324
rect 24737 1218 24771 1252
rect 24737 1146 24771 1180
rect 24737 1074 24771 1108
rect 24737 1002 24771 1036
rect 24867 1290 24901 1324
rect 24867 1218 24901 1252
rect 24867 1146 24901 1180
rect 24867 1074 24901 1108
rect 24867 1002 24901 1036
rect 24997 1290 25031 1324
rect 24997 1218 25031 1252
rect 24997 1146 25031 1180
rect 24997 1074 25031 1108
rect 24997 1002 25031 1036
rect 25127 1290 25161 1324
rect 25127 1218 25161 1252
rect 25127 1146 25161 1180
rect 25127 1074 25161 1108
rect 25127 1002 25161 1036
rect 25257 1290 25291 1324
rect 25257 1218 25291 1252
rect 25257 1146 25291 1180
rect 25257 1074 25291 1108
rect 25257 1002 25291 1036
rect 25387 1290 25421 1324
rect 25387 1218 25421 1252
rect 25387 1146 25421 1180
rect 25387 1074 25421 1108
rect 25387 1002 25421 1036
rect 25517 1290 25551 1324
rect 25517 1218 25551 1252
rect 25517 1146 25551 1180
rect 25517 1074 25551 1108
rect 25517 1002 25551 1036
rect 25647 1290 25681 1324
rect 25647 1218 25681 1252
rect 25647 1146 25681 1180
rect 25647 1074 25681 1108
rect 25647 1002 25681 1036
rect 25777 1290 25811 1324
rect 25777 1218 25811 1252
rect 25777 1146 25811 1180
rect 25777 1074 25811 1108
rect 25777 1002 25811 1036
rect 25907 1290 25941 1324
rect 25907 1218 25941 1252
rect 25907 1146 25941 1180
rect 25907 1074 25941 1108
rect 25907 1002 25941 1036
rect 26037 1290 26071 1324
rect 26037 1218 26071 1252
rect 26037 1146 26071 1180
rect 26037 1074 26071 1108
rect 26037 1002 26071 1036
rect 26167 1290 26201 1324
rect 26167 1218 26201 1252
rect 26167 1146 26201 1180
rect 26167 1074 26201 1108
rect 26167 1002 26201 1036
rect 26297 1290 26331 1324
rect 26297 1218 26331 1252
rect 26297 1146 26331 1180
rect 26297 1074 26331 1108
rect 26297 1002 26331 1036
rect 26427 1290 26461 1324
rect 26427 1218 26461 1252
rect 26427 1146 26461 1180
rect 26427 1074 26461 1108
rect 26427 1002 26461 1036
rect 26557 1290 26591 1324
rect 26557 1218 26591 1252
rect 26557 1146 26591 1180
rect 26557 1074 26591 1108
rect 26557 1002 26591 1036
rect 26687 1290 26721 1324
rect 26687 1218 26721 1252
rect 26687 1146 26721 1180
rect 26687 1074 26721 1108
rect 26687 1002 26721 1036
rect 26817 1290 26851 1324
rect 26817 1218 26851 1252
rect 26817 1146 26851 1180
rect 26817 1074 26851 1108
rect 26817 1002 26851 1036
rect 26947 1290 26981 1324
rect 26947 1218 26981 1252
rect 26947 1146 26981 1180
rect 26947 1074 26981 1108
rect 26947 1002 26981 1036
rect 27077 1290 27111 1324
rect 27077 1218 27111 1252
rect 27077 1146 27111 1180
rect 27077 1074 27111 1108
rect 27077 1002 27111 1036
rect 13210 873 13244 907
rect 13340 873 13374 907
rect 13470 873 13504 907
rect 13600 873 13634 907
rect 13730 873 13764 907
rect 13860 873 13894 907
rect 13990 873 14024 907
rect 14120 873 14154 907
rect 14250 873 14284 907
rect 14380 873 14414 907
rect 14510 873 14544 907
rect 14640 873 14674 907
rect 14770 873 14804 907
rect 14900 873 14934 907
rect 15030 873 15064 907
rect 15160 873 15194 907
rect 15290 873 15324 907
rect 15420 873 15454 907
rect 24802 873 24836 907
rect 24932 873 24966 907
rect 25062 873 25096 907
rect 25192 873 25226 907
rect 25322 873 25356 907
rect 25452 873 25486 907
rect 25582 873 25616 907
rect 25712 873 25746 907
rect 25842 873 25876 907
rect 25972 873 26006 907
rect 26102 873 26136 907
rect 26232 873 26266 907
rect 26362 873 26396 907
rect 26492 873 26526 907
rect 26622 873 26656 907
rect 26752 873 26786 907
rect 26882 873 26916 907
rect 27012 873 27046 907
rect 13196 740 13204 774
rect 13204 740 13230 774
rect 13268 740 13272 774
rect 13272 740 13302 774
rect 13340 740 13374 774
rect 13412 740 13442 774
rect 13442 740 13446 774
rect 13484 740 13510 774
rect 13510 740 13518 774
rect 13586 740 13594 774
rect 13594 740 13620 774
rect 13658 740 13662 774
rect 13662 740 13692 774
rect 13730 740 13764 774
rect 13802 740 13832 774
rect 13832 740 13836 774
rect 13874 740 13900 774
rect 13900 740 13908 774
rect 13976 740 13984 774
rect 13984 740 14010 774
rect 14048 740 14052 774
rect 14052 740 14082 774
rect 14120 740 14154 774
rect 14192 740 14222 774
rect 14222 740 14226 774
rect 14264 740 14290 774
rect 14290 740 14298 774
rect 14366 740 14374 774
rect 14374 740 14400 774
rect 14438 740 14442 774
rect 14442 740 14472 774
rect 14510 740 14544 774
rect 14582 740 14612 774
rect 14612 740 14616 774
rect 14654 740 14680 774
rect 14680 740 14688 774
rect 14756 740 14764 774
rect 14764 740 14790 774
rect 14828 740 14832 774
rect 14832 740 14862 774
rect 14900 740 14934 774
rect 14972 740 15002 774
rect 15002 740 15006 774
rect 15044 740 15070 774
rect 15070 740 15078 774
rect 15146 740 15154 774
rect 15154 740 15180 774
rect 15218 740 15222 774
rect 15222 740 15252 774
rect 15290 740 15324 774
rect 15362 740 15392 774
rect 15392 740 15396 774
rect 15434 740 15460 774
rect 15460 740 15468 774
rect 24788 740 24796 774
rect 24796 740 24822 774
rect 24860 740 24864 774
rect 24864 740 24894 774
rect 24932 740 24966 774
rect 25004 740 25034 774
rect 25034 740 25038 774
rect 25076 740 25102 774
rect 25102 740 25110 774
rect 25178 740 25186 774
rect 25186 740 25212 774
rect 25250 740 25254 774
rect 25254 740 25284 774
rect 25322 740 25356 774
rect 25394 740 25424 774
rect 25424 740 25428 774
rect 25466 740 25492 774
rect 25492 740 25500 774
rect 25568 740 25576 774
rect 25576 740 25602 774
rect 25640 740 25644 774
rect 25644 740 25674 774
rect 25712 740 25746 774
rect 25784 740 25814 774
rect 25814 740 25818 774
rect 25856 740 25882 774
rect 25882 740 25890 774
rect 25958 740 25966 774
rect 25966 740 25992 774
rect 26030 740 26034 774
rect 26034 740 26064 774
rect 26102 740 26136 774
rect 26174 740 26204 774
rect 26204 740 26208 774
rect 26246 740 26272 774
rect 26272 740 26280 774
rect 26348 740 26356 774
rect 26356 740 26382 774
rect 26420 740 26424 774
rect 26424 740 26454 774
rect 26492 740 26526 774
rect 26564 740 26594 774
rect 26594 740 26598 774
rect 26636 740 26662 774
rect 26662 740 26670 774
rect 26738 740 26746 774
rect 26746 740 26772 774
rect 26810 740 26814 774
rect 26814 740 26844 774
rect 26882 740 26916 774
rect 26954 740 26984 774
rect 26984 740 26988 774
rect 27026 740 27052 774
rect 27052 740 27060 774
<< metal1 >>
rect 12823 5495 15593 5509
rect 12823 5443 12833 5495
rect 12885 5443 12897 5495
rect 12949 5443 12961 5495
rect 13013 5486 13657 5495
rect 13013 5452 13022 5486
rect 13056 5452 13104 5486
rect 13138 5452 13196 5486
rect 13230 5452 13268 5486
rect 13302 5452 13340 5486
rect 13374 5452 13412 5486
rect 13446 5452 13484 5486
rect 13518 5452 13586 5486
rect 13620 5452 13657 5486
rect 13013 5443 13657 5452
rect 13709 5443 13721 5495
rect 13773 5443 13785 5495
rect 13837 5486 14437 5495
rect 13837 5452 13874 5486
rect 13908 5452 13976 5486
rect 14010 5452 14048 5486
rect 14082 5452 14120 5486
rect 14154 5452 14192 5486
rect 14226 5452 14264 5486
rect 14298 5452 14366 5486
rect 14400 5452 14437 5486
rect 13837 5443 14437 5452
rect 14489 5443 14501 5495
rect 14553 5443 14565 5495
rect 14617 5486 15217 5495
rect 14617 5452 14654 5486
rect 14688 5452 14756 5486
rect 14790 5452 14828 5486
rect 14862 5452 14900 5486
rect 14934 5452 14972 5486
rect 15006 5452 15044 5486
rect 15078 5452 15217 5486
rect 14617 5443 15217 5452
rect 15269 5443 15281 5495
rect 15333 5443 15345 5495
rect 15397 5443 15593 5495
rect 12823 5429 15593 5443
rect 24415 5495 27185 5509
rect 24415 5443 24425 5495
rect 24477 5443 24489 5495
rect 24541 5443 24553 5495
rect 24605 5486 25249 5495
rect 24605 5452 24614 5486
rect 24648 5452 24696 5486
rect 24730 5452 24788 5486
rect 24822 5452 24860 5486
rect 24894 5452 24932 5486
rect 24966 5452 25004 5486
rect 25038 5452 25076 5486
rect 25110 5452 25178 5486
rect 25212 5452 25249 5486
rect 24605 5443 25249 5452
rect 25301 5443 25313 5495
rect 25365 5443 25377 5495
rect 25429 5486 26029 5495
rect 25429 5452 25466 5486
rect 25500 5452 25568 5486
rect 25602 5452 25640 5486
rect 25674 5452 25712 5486
rect 25746 5452 25784 5486
rect 25818 5452 25856 5486
rect 25890 5452 25958 5486
rect 25992 5452 26029 5486
rect 25429 5443 26029 5452
rect 26081 5443 26093 5495
rect 26145 5443 26157 5495
rect 26209 5486 26809 5495
rect 26209 5452 26246 5486
rect 26280 5452 26348 5486
rect 26382 5452 26420 5486
rect 26454 5452 26492 5486
rect 26526 5452 26564 5486
rect 26598 5452 26636 5486
rect 26670 5452 26809 5486
rect 26209 5443 26809 5452
rect 26861 5443 26873 5495
rect 26925 5443 26937 5495
rect 26989 5443 27185 5495
rect 24415 5429 27185 5443
rect 12493 5362 12567 5369
rect 12493 5310 12504 5362
rect 12556 5310 12567 5362
rect 12493 5303 12567 5310
rect 13000 5362 13134 5369
rect 13000 5310 13009 5362
rect 13061 5310 13073 5362
rect 13125 5310 13134 5362
rect 13190 5353 13264 5429
rect 13190 5319 13210 5353
rect 13244 5319 13264 5353
rect 13190 5313 13264 5319
rect 13320 5362 13394 5369
rect 13000 5303 13134 5310
rect 13320 5310 13331 5362
rect 13383 5310 13394 5362
rect 13450 5353 13524 5429
rect 13450 5319 13470 5353
rect 13504 5319 13524 5353
rect 13450 5313 13524 5319
rect 13580 5353 13654 5429
rect 13580 5319 13600 5353
rect 13634 5319 13654 5353
rect 13580 5313 13654 5319
rect 13710 5362 13784 5369
rect 13320 5303 13394 5310
rect 13710 5310 13721 5362
rect 13773 5310 13784 5362
rect 13840 5353 13914 5429
rect 13840 5319 13860 5353
rect 13894 5319 13914 5353
rect 13840 5313 13914 5319
rect 13970 5353 14044 5429
rect 13970 5319 13990 5353
rect 14024 5319 14044 5353
rect 13970 5313 14044 5319
rect 14100 5362 14174 5369
rect 13710 5303 13784 5310
rect 14100 5310 14111 5362
rect 14163 5310 14174 5362
rect 14230 5353 14304 5429
rect 14230 5319 14250 5353
rect 14284 5319 14304 5353
rect 14230 5313 14304 5319
rect 14360 5353 14434 5429
rect 14360 5319 14380 5353
rect 14414 5319 14434 5353
rect 14360 5313 14434 5319
rect 14490 5362 14564 5369
rect 14100 5303 14174 5310
rect 14490 5310 14501 5362
rect 14553 5310 14564 5362
rect 14620 5353 14694 5429
rect 14620 5319 14640 5353
rect 14674 5319 14694 5353
rect 14620 5313 14694 5319
rect 14750 5353 14824 5429
rect 14750 5319 14770 5353
rect 14804 5319 14824 5353
rect 14750 5313 14824 5319
rect 14880 5362 14954 5369
rect 14490 5303 14564 5310
rect 14880 5310 14891 5362
rect 14943 5310 14954 5362
rect 15010 5353 15084 5429
rect 15010 5319 15030 5353
rect 15064 5319 15084 5353
rect 15010 5313 15084 5319
rect 24085 5362 24159 5369
rect 14880 5303 14954 5310
rect 24085 5310 24096 5362
rect 24148 5310 24159 5362
rect 24085 5303 24159 5310
rect 24592 5362 24726 5369
rect 24592 5310 24601 5362
rect 24653 5310 24665 5362
rect 24717 5310 24726 5362
rect 24782 5353 24856 5429
rect 24782 5319 24802 5353
rect 24836 5319 24856 5353
rect 24782 5313 24856 5319
rect 24912 5362 24986 5369
rect 24592 5303 24726 5310
rect 24912 5310 24923 5362
rect 24975 5310 24986 5362
rect 25042 5353 25116 5429
rect 25042 5319 25062 5353
rect 25096 5319 25116 5353
rect 25042 5313 25116 5319
rect 25172 5353 25246 5429
rect 25172 5319 25192 5353
rect 25226 5319 25246 5353
rect 25172 5313 25246 5319
rect 25302 5362 25376 5369
rect 24912 5303 24986 5310
rect 25302 5310 25313 5362
rect 25365 5310 25376 5362
rect 25432 5353 25506 5429
rect 25432 5319 25452 5353
rect 25486 5319 25506 5353
rect 25432 5313 25506 5319
rect 25562 5353 25636 5429
rect 25562 5319 25582 5353
rect 25616 5319 25636 5353
rect 25562 5313 25636 5319
rect 25692 5362 25766 5369
rect 25302 5303 25376 5310
rect 25692 5310 25703 5362
rect 25755 5310 25766 5362
rect 25822 5353 25896 5429
rect 25822 5319 25842 5353
rect 25876 5319 25896 5353
rect 25822 5313 25896 5319
rect 25952 5353 26026 5429
rect 25952 5319 25972 5353
rect 26006 5319 26026 5353
rect 25952 5313 26026 5319
rect 26082 5362 26156 5369
rect 25692 5303 25766 5310
rect 26082 5310 26093 5362
rect 26145 5310 26156 5362
rect 26212 5353 26286 5429
rect 26212 5319 26232 5353
rect 26266 5319 26286 5353
rect 26212 5313 26286 5319
rect 26342 5353 26416 5429
rect 26342 5319 26362 5353
rect 26396 5319 26416 5353
rect 26342 5313 26416 5319
rect 26472 5362 26546 5369
rect 26082 5303 26156 5310
rect 26472 5310 26483 5362
rect 26535 5310 26546 5362
rect 26602 5353 26676 5429
rect 26602 5319 26622 5353
rect 26656 5319 26676 5353
rect 26602 5313 26676 5319
rect 26472 5303 26546 5310
rect 13000 5224 13064 5236
rect 13000 5217 13015 5224
rect 13049 5217 13064 5224
rect 13000 5165 13006 5217
rect 13058 5165 13064 5217
rect 13000 5153 13064 5165
rect 13000 5101 13006 5153
rect 13058 5101 13064 5153
rect 13139 5224 13185 5236
rect 13139 5190 13145 5224
rect 13179 5190 13185 5224
rect 13139 5152 13185 5190
rect 13139 5118 13145 5152
rect 13179 5118 13185 5152
rect 13139 5113 13185 5118
rect 13269 5224 13315 5236
rect 13269 5190 13275 5224
rect 13309 5190 13315 5224
rect 13269 5152 13315 5190
rect 13269 5118 13275 5152
rect 13309 5118 13315 5152
rect 13000 5089 13064 5101
rect 13000 5037 13006 5089
rect 13058 5037 13064 5089
rect 13000 5025 13064 5037
rect 13000 4973 13006 5025
rect 13058 4973 13064 5025
rect 13125 5089 13199 5113
rect 13125 5037 13136 5089
rect 13188 5037 13199 5089
rect 13125 5013 13199 5037
rect 13269 5080 13315 5118
rect 13399 5224 13445 5236
rect 13399 5190 13405 5224
rect 13439 5190 13445 5224
rect 13399 5152 13445 5190
rect 13399 5118 13405 5152
rect 13439 5118 13445 5152
rect 13399 5113 13445 5118
rect 13529 5224 13575 5236
rect 13529 5190 13535 5224
rect 13569 5190 13575 5224
rect 13529 5152 13575 5190
rect 13529 5118 13535 5152
rect 13569 5118 13575 5152
rect 13529 5113 13575 5118
rect 13659 5224 13705 5236
rect 13659 5190 13665 5224
rect 13699 5190 13705 5224
rect 13659 5152 13705 5190
rect 13659 5118 13665 5152
rect 13699 5118 13705 5152
rect 13269 5046 13275 5080
rect 13309 5046 13315 5080
rect 13000 4961 13064 4973
rect 13000 4909 13006 4961
rect 13058 4909 13064 4961
rect 13000 4902 13015 4909
rect 13049 4902 13064 4909
rect 13000 4890 13064 4902
rect 13139 5008 13185 5013
rect 13139 4974 13145 5008
rect 13179 4974 13185 5008
rect 13139 4936 13185 4974
rect 13139 4902 13145 4936
rect 13179 4902 13185 4936
rect 13139 4890 13185 4902
rect 13269 5008 13315 5046
rect 13385 5089 13459 5113
rect 13385 5037 13396 5089
rect 13448 5037 13459 5089
rect 13385 5013 13459 5037
rect 13515 5089 13589 5113
rect 13515 5037 13526 5089
rect 13578 5037 13589 5089
rect 13515 5013 13589 5037
rect 13659 5080 13705 5118
rect 13789 5224 13835 5236
rect 13789 5190 13795 5224
rect 13829 5190 13835 5224
rect 13789 5152 13835 5190
rect 13789 5118 13795 5152
rect 13829 5118 13835 5152
rect 13789 5113 13835 5118
rect 13919 5224 13965 5236
rect 13919 5190 13925 5224
rect 13959 5190 13965 5224
rect 13919 5152 13965 5190
rect 13919 5118 13925 5152
rect 13959 5118 13965 5152
rect 13919 5113 13965 5118
rect 14049 5224 14095 5236
rect 14049 5190 14055 5224
rect 14089 5190 14095 5224
rect 14049 5152 14095 5190
rect 14049 5118 14055 5152
rect 14089 5118 14095 5152
rect 13659 5046 13665 5080
rect 13699 5046 13705 5080
rect 13269 4974 13275 5008
rect 13309 4974 13315 5008
rect 13269 4936 13315 4974
rect 13269 4902 13275 4936
rect 13309 4902 13315 4936
rect 13269 4676 13315 4902
rect 13399 5008 13445 5013
rect 13399 4974 13405 5008
rect 13439 4974 13445 5008
rect 13399 4936 13445 4974
rect 13399 4902 13405 4936
rect 13439 4902 13445 4936
rect 13399 4890 13445 4902
rect 13529 5008 13575 5013
rect 13529 4974 13535 5008
rect 13569 4974 13575 5008
rect 13529 4936 13575 4974
rect 13529 4902 13535 4936
rect 13569 4902 13575 4936
rect 13529 4890 13575 4902
rect 13659 5008 13705 5046
rect 13775 5089 13849 5113
rect 13775 5037 13786 5089
rect 13838 5037 13849 5089
rect 13775 5013 13849 5037
rect 13905 5089 13979 5113
rect 13905 5037 13916 5089
rect 13968 5037 13979 5089
rect 13905 5013 13979 5037
rect 14049 5080 14095 5118
rect 14179 5224 14225 5236
rect 14179 5190 14185 5224
rect 14219 5190 14225 5224
rect 14179 5152 14225 5190
rect 14179 5118 14185 5152
rect 14219 5118 14225 5152
rect 14179 5113 14225 5118
rect 14309 5224 14355 5236
rect 14309 5190 14315 5224
rect 14349 5190 14355 5224
rect 14309 5152 14355 5190
rect 14309 5118 14315 5152
rect 14349 5118 14355 5152
rect 14309 5113 14355 5118
rect 14439 5224 14485 5236
rect 14439 5190 14445 5224
rect 14479 5190 14485 5224
rect 14439 5152 14485 5190
rect 14439 5118 14445 5152
rect 14479 5118 14485 5152
rect 14049 5046 14055 5080
rect 14089 5046 14095 5080
rect 13659 4974 13665 5008
rect 13699 4974 13705 5008
rect 13659 4936 13705 4974
rect 13659 4902 13665 4936
rect 13699 4902 13705 4936
rect 13269 4642 13275 4676
rect 13309 4642 13315 4676
rect 13269 4604 13315 4642
rect 13269 4570 13275 4604
rect 13309 4570 13315 4604
rect 13269 4532 13315 4570
rect 13269 4498 13275 4532
rect 13309 4498 13315 4532
rect 13269 4460 13315 4498
rect 13269 4426 13275 4460
rect 13309 4426 13315 4460
rect 13269 4388 13315 4426
rect 13269 4354 13275 4388
rect 13309 4354 13315 4388
rect 13269 4342 13315 4354
rect 13390 4676 13454 4688
rect 13390 4669 13405 4676
rect 13439 4669 13454 4676
rect 13390 4617 13396 4669
rect 13448 4617 13454 4669
rect 13390 4605 13454 4617
rect 13390 4553 13396 4605
rect 13448 4553 13454 4605
rect 13390 4541 13454 4553
rect 13390 4489 13396 4541
rect 13448 4489 13454 4541
rect 13390 4477 13454 4489
rect 13390 4425 13396 4477
rect 13448 4425 13454 4477
rect 13390 4413 13454 4425
rect 13390 4361 13396 4413
rect 13448 4361 13454 4413
rect 13390 4354 13405 4361
rect 13439 4354 13454 4361
rect 13390 4342 13454 4354
rect 13659 4676 13705 4902
rect 13789 5008 13835 5013
rect 13789 4974 13795 5008
rect 13829 4974 13835 5008
rect 13789 4936 13835 4974
rect 13789 4902 13795 4936
rect 13829 4902 13835 4936
rect 13789 4890 13835 4902
rect 13919 5008 13965 5013
rect 13919 4974 13925 5008
rect 13959 4974 13965 5008
rect 13919 4936 13965 4974
rect 13919 4902 13925 4936
rect 13959 4902 13965 4936
rect 13919 4890 13965 4902
rect 14049 5008 14095 5046
rect 14165 5089 14239 5113
rect 14165 5037 14176 5089
rect 14228 5037 14239 5089
rect 14165 5013 14239 5037
rect 14295 5089 14369 5113
rect 14295 5037 14306 5089
rect 14358 5037 14369 5089
rect 14295 5013 14369 5037
rect 14439 5080 14485 5118
rect 14569 5224 14615 5236
rect 14569 5190 14575 5224
rect 14609 5190 14615 5224
rect 14569 5152 14615 5190
rect 14569 5118 14575 5152
rect 14609 5118 14615 5152
rect 14569 5113 14615 5118
rect 14699 5224 14745 5236
rect 14699 5190 14705 5224
rect 14739 5190 14745 5224
rect 14699 5152 14745 5190
rect 14699 5118 14705 5152
rect 14739 5118 14745 5152
rect 14699 5113 14745 5118
rect 14829 5224 14875 5236
rect 14829 5190 14835 5224
rect 14869 5190 14875 5224
rect 14829 5152 14875 5190
rect 14829 5118 14835 5152
rect 14869 5118 14875 5152
rect 14439 5046 14445 5080
rect 14479 5046 14485 5080
rect 14049 4974 14055 5008
rect 14089 4974 14095 5008
rect 14049 4936 14095 4974
rect 14049 4902 14055 4936
rect 14089 4902 14095 4936
rect 13659 4642 13665 4676
rect 13699 4642 13705 4676
rect 13659 4604 13705 4642
rect 13659 4570 13665 4604
rect 13699 4570 13705 4604
rect 13659 4532 13705 4570
rect 13659 4498 13665 4532
rect 13699 4498 13705 4532
rect 13659 4460 13705 4498
rect 13659 4426 13665 4460
rect 13699 4426 13705 4460
rect 13659 4388 13705 4426
rect 13659 4354 13665 4388
rect 13699 4354 13705 4388
rect 13659 4342 13705 4354
rect 13780 4676 13844 4688
rect 13780 4669 13795 4676
rect 13829 4669 13844 4676
rect 13780 4617 13786 4669
rect 13838 4617 13844 4669
rect 13780 4605 13844 4617
rect 13780 4553 13786 4605
rect 13838 4553 13844 4605
rect 13780 4541 13844 4553
rect 13780 4489 13786 4541
rect 13838 4489 13844 4541
rect 13780 4477 13844 4489
rect 13780 4425 13786 4477
rect 13838 4425 13844 4477
rect 13780 4413 13844 4425
rect 13780 4361 13786 4413
rect 13838 4361 13844 4413
rect 13780 4354 13795 4361
rect 13829 4354 13844 4361
rect 13780 4342 13844 4354
rect 14049 4676 14095 4902
rect 14179 5008 14225 5013
rect 14179 4974 14185 5008
rect 14219 4974 14225 5008
rect 14179 4936 14225 4974
rect 14179 4902 14185 4936
rect 14219 4902 14225 4936
rect 14179 4890 14225 4902
rect 14309 5008 14355 5013
rect 14309 4974 14315 5008
rect 14349 4974 14355 5008
rect 14309 4936 14355 4974
rect 14309 4902 14315 4936
rect 14349 4902 14355 4936
rect 14309 4890 14355 4902
rect 14439 5008 14485 5046
rect 14555 5089 14629 5113
rect 14555 5037 14566 5089
rect 14618 5037 14629 5089
rect 14555 5013 14629 5037
rect 14685 5089 14759 5113
rect 14685 5037 14696 5089
rect 14748 5037 14759 5089
rect 14685 5013 14759 5037
rect 14829 5080 14875 5118
rect 14959 5224 15005 5236
rect 14959 5190 14965 5224
rect 14999 5190 15005 5224
rect 14959 5152 15005 5190
rect 14959 5118 14965 5152
rect 14999 5118 15005 5152
rect 14959 5113 15005 5118
rect 15089 5224 15135 5236
rect 15089 5190 15095 5224
rect 15129 5190 15135 5224
rect 15089 5152 15135 5190
rect 15089 5118 15095 5152
rect 15129 5118 15135 5152
rect 15089 5113 15135 5118
rect 24592 5224 24656 5236
rect 24592 5217 24607 5224
rect 24641 5217 24656 5224
rect 24592 5165 24598 5217
rect 24650 5165 24656 5217
rect 24592 5153 24656 5165
rect 14829 5046 14835 5080
rect 14869 5046 14875 5080
rect 14439 4974 14445 5008
rect 14479 4974 14485 5008
rect 14439 4936 14485 4974
rect 14439 4902 14445 4936
rect 14479 4902 14485 4936
rect 14049 4642 14055 4676
rect 14089 4642 14095 4676
rect 14049 4604 14095 4642
rect 14049 4570 14055 4604
rect 14089 4570 14095 4604
rect 14049 4532 14095 4570
rect 14049 4498 14055 4532
rect 14089 4498 14095 4532
rect 14049 4460 14095 4498
rect 14049 4426 14055 4460
rect 14089 4426 14095 4460
rect 14049 4388 14095 4426
rect 14049 4354 14055 4388
rect 14089 4354 14095 4388
rect 14049 4342 14095 4354
rect 14170 4676 14234 4688
rect 14170 4669 14185 4676
rect 14219 4669 14234 4676
rect 14170 4617 14176 4669
rect 14228 4617 14234 4669
rect 14170 4605 14234 4617
rect 14170 4553 14176 4605
rect 14228 4553 14234 4605
rect 14170 4541 14234 4553
rect 14170 4489 14176 4541
rect 14228 4489 14234 4541
rect 14170 4477 14234 4489
rect 14170 4425 14176 4477
rect 14228 4425 14234 4477
rect 14170 4413 14234 4425
rect 14170 4361 14176 4413
rect 14228 4361 14234 4413
rect 14170 4354 14185 4361
rect 14219 4354 14234 4361
rect 14170 4342 14234 4354
rect 14439 4676 14485 4902
rect 14569 5008 14615 5013
rect 14569 4974 14575 5008
rect 14609 4974 14615 5008
rect 14569 4936 14615 4974
rect 14569 4902 14575 4936
rect 14609 4902 14615 4936
rect 14569 4890 14615 4902
rect 14699 5008 14745 5013
rect 14699 4974 14705 5008
rect 14739 4974 14745 5008
rect 14699 4936 14745 4974
rect 14699 4902 14705 4936
rect 14739 4902 14745 4936
rect 14699 4890 14745 4902
rect 14829 5008 14875 5046
rect 14945 5089 15019 5113
rect 14945 5037 14956 5089
rect 15008 5037 15019 5089
rect 14945 5013 15019 5037
rect 15075 5089 15149 5113
rect 15075 5037 15086 5089
rect 15138 5037 15149 5089
rect 15075 5013 15149 5037
rect 24592 5101 24598 5153
rect 24650 5101 24656 5153
rect 24731 5224 24777 5236
rect 24731 5190 24737 5224
rect 24771 5190 24777 5224
rect 24731 5152 24777 5190
rect 24731 5118 24737 5152
rect 24771 5118 24777 5152
rect 24731 5113 24777 5118
rect 24861 5224 24907 5236
rect 24861 5190 24867 5224
rect 24901 5190 24907 5224
rect 24861 5152 24907 5190
rect 24861 5118 24867 5152
rect 24901 5118 24907 5152
rect 24592 5089 24656 5101
rect 24592 5037 24598 5089
rect 24650 5037 24656 5089
rect 24592 5025 24656 5037
rect 14829 4974 14835 5008
rect 14869 4974 14875 5008
rect 14829 4936 14875 4974
rect 14829 4902 14835 4936
rect 14869 4902 14875 4936
rect 14439 4642 14445 4676
rect 14479 4642 14485 4676
rect 14439 4604 14485 4642
rect 14439 4570 14445 4604
rect 14479 4570 14485 4604
rect 14439 4532 14485 4570
rect 14439 4498 14445 4532
rect 14479 4498 14485 4532
rect 14439 4460 14485 4498
rect 14439 4426 14445 4460
rect 14479 4426 14485 4460
rect 14439 4388 14485 4426
rect 14439 4354 14445 4388
rect 14479 4354 14485 4388
rect 14439 4342 14485 4354
rect 14560 4676 14624 4688
rect 14560 4669 14575 4676
rect 14609 4669 14624 4676
rect 14560 4617 14566 4669
rect 14618 4617 14624 4669
rect 14560 4605 14624 4617
rect 14560 4553 14566 4605
rect 14618 4553 14624 4605
rect 14560 4541 14624 4553
rect 14560 4489 14566 4541
rect 14618 4489 14624 4541
rect 14560 4477 14624 4489
rect 14560 4425 14566 4477
rect 14618 4425 14624 4477
rect 14560 4413 14624 4425
rect 14560 4361 14566 4413
rect 14618 4361 14624 4413
rect 14560 4354 14575 4361
rect 14609 4354 14624 4361
rect 14560 4342 14624 4354
rect 14829 4676 14875 4902
rect 14959 5008 15005 5013
rect 14959 4974 14965 5008
rect 14999 4974 15005 5008
rect 14959 4936 15005 4974
rect 14959 4902 14965 4936
rect 14999 4902 15005 4936
rect 14959 4890 15005 4902
rect 15089 5008 15135 5013
rect 15089 4974 15095 5008
rect 15129 4974 15135 5008
rect 15089 4936 15135 4974
rect 15089 4902 15095 4936
rect 15129 4902 15135 4936
rect 24592 4973 24598 5025
rect 24650 4973 24656 5025
rect 24717 5089 24791 5113
rect 24717 5037 24728 5089
rect 24780 5037 24791 5089
rect 24717 5013 24791 5037
rect 24861 5080 24907 5118
rect 24991 5224 25037 5236
rect 24991 5190 24997 5224
rect 25031 5190 25037 5224
rect 24991 5152 25037 5190
rect 24991 5118 24997 5152
rect 25031 5118 25037 5152
rect 24991 5113 25037 5118
rect 25121 5224 25167 5236
rect 25121 5190 25127 5224
rect 25161 5190 25167 5224
rect 25121 5152 25167 5190
rect 25121 5118 25127 5152
rect 25161 5118 25167 5152
rect 25121 5113 25167 5118
rect 25251 5224 25297 5236
rect 25251 5190 25257 5224
rect 25291 5190 25297 5224
rect 25251 5152 25297 5190
rect 25251 5118 25257 5152
rect 25291 5118 25297 5152
rect 24861 5046 24867 5080
rect 24901 5046 24907 5080
rect 24592 4961 24656 4973
rect 15089 4890 15135 4902
rect 15284 4924 15524 4927
rect 15284 4915 15317 4924
rect 15284 4881 15315 4915
rect 15284 4872 15317 4881
rect 15369 4872 15381 4924
rect 15433 4872 15445 4924
rect 15497 4872 15524 4924
rect 24592 4909 24598 4961
rect 24650 4909 24656 4961
rect 24592 4902 24607 4909
rect 24641 4902 24656 4909
rect 24592 4890 24656 4902
rect 24731 5008 24777 5013
rect 24731 4974 24737 5008
rect 24771 4974 24777 5008
rect 24731 4936 24777 4974
rect 24731 4902 24737 4936
rect 24771 4902 24777 4936
rect 24731 4890 24777 4902
rect 24861 5008 24907 5046
rect 24977 5089 25051 5113
rect 24977 5037 24988 5089
rect 25040 5037 25051 5089
rect 24977 5013 25051 5037
rect 25107 5089 25181 5113
rect 25107 5037 25118 5089
rect 25170 5037 25181 5089
rect 25107 5013 25181 5037
rect 25251 5080 25297 5118
rect 25381 5224 25427 5236
rect 25381 5190 25387 5224
rect 25421 5190 25427 5224
rect 25381 5152 25427 5190
rect 25381 5118 25387 5152
rect 25421 5118 25427 5152
rect 25381 5113 25427 5118
rect 25511 5224 25557 5236
rect 25511 5190 25517 5224
rect 25551 5190 25557 5224
rect 25511 5152 25557 5190
rect 25511 5118 25517 5152
rect 25551 5118 25557 5152
rect 25511 5113 25557 5118
rect 25641 5224 25687 5236
rect 25641 5190 25647 5224
rect 25681 5190 25687 5224
rect 25641 5152 25687 5190
rect 25641 5118 25647 5152
rect 25681 5118 25687 5152
rect 25251 5046 25257 5080
rect 25291 5046 25297 5080
rect 24861 4974 24867 5008
rect 24901 4974 24907 5008
rect 24861 4936 24907 4974
rect 24861 4902 24867 4936
rect 24901 4902 24907 4936
rect 15284 4869 15524 4872
rect 15198 4781 15204 4833
rect 15256 4827 15262 4833
rect 15375 4827 15535 4834
rect 15256 4824 15535 4827
rect 15256 4790 15402 4824
rect 15436 4790 15474 4824
rect 15508 4790 15535 4824
rect 15256 4787 15535 4790
rect 15256 4781 15262 4787
rect 15375 4780 15535 4787
rect 14829 4642 14835 4676
rect 14869 4642 14875 4676
rect 14829 4604 14875 4642
rect 14829 4570 14835 4604
rect 14869 4570 14875 4604
rect 14829 4532 14875 4570
rect 14829 4498 14835 4532
rect 14869 4498 14875 4532
rect 14829 4460 14875 4498
rect 14829 4426 14835 4460
rect 14869 4426 14875 4460
rect 14829 4388 14875 4426
rect 14829 4354 14835 4388
rect 14869 4354 14875 4388
rect 14829 4342 14875 4354
rect 14950 4676 15014 4688
rect 14950 4669 14965 4676
rect 14999 4669 15014 4676
rect 14950 4617 14956 4669
rect 15008 4617 15014 4669
rect 14950 4605 15014 4617
rect 14950 4553 14956 4605
rect 15008 4553 15014 4605
rect 14950 4541 15014 4553
rect 14950 4489 14956 4541
rect 15008 4489 15014 4541
rect 14950 4477 15014 4489
rect 14950 4425 14956 4477
rect 15008 4425 15014 4477
rect 14950 4413 15014 4425
rect 14950 4361 14956 4413
rect 15008 4361 15014 4413
rect 15203 4676 15249 4688
rect 15293 4685 15339 4688
rect 15203 4642 15209 4676
rect 15243 4642 15249 4676
rect 15203 4604 15249 4642
rect 15284 4633 15290 4685
rect 15342 4633 15348 4685
rect 15383 4676 15429 4688
rect 15473 4685 15519 4688
rect 15383 4642 15389 4676
rect 15423 4642 15429 4676
rect 15203 4570 15209 4604
rect 15243 4570 15249 4604
rect 15203 4532 15249 4570
rect 15203 4498 15209 4532
rect 15243 4498 15249 4532
rect 15203 4460 15249 4498
rect 15203 4426 15209 4460
rect 15243 4426 15249 4460
rect 15203 4397 15249 4426
rect 15293 4604 15339 4633
rect 15293 4570 15299 4604
rect 15333 4570 15339 4604
rect 15293 4532 15339 4570
rect 15293 4498 15299 4532
rect 15333 4498 15339 4532
rect 15293 4460 15339 4498
rect 15293 4426 15299 4460
rect 15333 4426 15339 4460
rect 14950 4354 14965 4361
rect 14999 4354 15014 4361
rect 14950 4342 15014 4354
rect 15194 4345 15200 4397
rect 15252 4345 15258 4397
rect 15293 4388 15339 4426
rect 15383 4604 15429 4642
rect 15464 4633 15470 4685
rect 15522 4633 15528 4685
rect 15563 4676 15609 4688
rect 15563 4642 15569 4676
rect 15603 4642 15609 4676
rect 15383 4570 15389 4604
rect 15423 4570 15429 4604
rect 15383 4532 15429 4570
rect 15383 4498 15389 4532
rect 15423 4498 15429 4532
rect 15383 4460 15429 4498
rect 15383 4426 15389 4460
rect 15423 4426 15429 4460
rect 15383 4392 15429 4426
rect 15473 4604 15519 4633
rect 15473 4570 15479 4604
rect 15513 4570 15519 4604
rect 15473 4532 15519 4570
rect 15473 4498 15479 4532
rect 15513 4498 15519 4532
rect 15473 4460 15519 4498
rect 15473 4426 15479 4460
rect 15513 4426 15519 4460
rect 15293 4354 15299 4388
rect 15333 4354 15339 4388
rect 15203 4342 15249 4345
rect 15293 4342 15339 4354
rect 15373 4391 15439 4392
rect 15373 4339 15380 4391
rect 15432 4339 15439 4391
rect 15473 4388 15519 4426
rect 15563 4604 15609 4642
rect 15563 4570 15569 4604
rect 15603 4570 15609 4604
rect 15563 4532 15609 4570
rect 15563 4498 15569 4532
rect 15603 4498 15609 4532
rect 15563 4460 15609 4498
rect 15563 4426 15569 4460
rect 15603 4426 15609 4460
rect 15563 4392 15609 4426
rect 24861 4676 24907 4902
rect 24991 5008 25037 5013
rect 24991 4974 24997 5008
rect 25031 4974 25037 5008
rect 24991 4936 25037 4974
rect 24991 4902 24997 4936
rect 25031 4902 25037 4936
rect 24991 4890 25037 4902
rect 25121 5008 25167 5013
rect 25121 4974 25127 5008
rect 25161 4974 25167 5008
rect 25121 4936 25167 4974
rect 25121 4902 25127 4936
rect 25161 4902 25167 4936
rect 25121 4890 25167 4902
rect 25251 5008 25297 5046
rect 25367 5089 25441 5113
rect 25367 5037 25378 5089
rect 25430 5037 25441 5089
rect 25367 5013 25441 5037
rect 25497 5089 25571 5113
rect 25497 5037 25508 5089
rect 25560 5037 25571 5089
rect 25497 5013 25571 5037
rect 25641 5080 25687 5118
rect 25771 5224 25817 5236
rect 25771 5190 25777 5224
rect 25811 5190 25817 5224
rect 25771 5152 25817 5190
rect 25771 5118 25777 5152
rect 25811 5118 25817 5152
rect 25771 5113 25817 5118
rect 25901 5224 25947 5236
rect 25901 5190 25907 5224
rect 25941 5190 25947 5224
rect 25901 5152 25947 5190
rect 25901 5118 25907 5152
rect 25941 5118 25947 5152
rect 25901 5113 25947 5118
rect 26031 5224 26077 5236
rect 26031 5190 26037 5224
rect 26071 5190 26077 5224
rect 26031 5152 26077 5190
rect 26031 5118 26037 5152
rect 26071 5118 26077 5152
rect 25641 5046 25647 5080
rect 25681 5046 25687 5080
rect 25251 4974 25257 5008
rect 25291 4974 25297 5008
rect 25251 4936 25297 4974
rect 25251 4902 25257 4936
rect 25291 4902 25297 4936
rect 24861 4642 24867 4676
rect 24901 4642 24907 4676
rect 24861 4604 24907 4642
rect 24861 4570 24867 4604
rect 24901 4570 24907 4604
rect 24861 4532 24907 4570
rect 24861 4498 24867 4532
rect 24901 4498 24907 4532
rect 24861 4460 24907 4498
rect 24861 4426 24867 4460
rect 24901 4426 24907 4460
rect 15473 4354 15479 4388
rect 15513 4354 15519 4388
rect 15473 4342 15519 4354
rect 15553 4391 15619 4392
rect 15373 4338 15439 4339
rect 15553 4339 15560 4391
rect 15612 4339 15619 4391
rect 24861 4388 24907 4426
rect 24861 4354 24867 4388
rect 24901 4354 24907 4388
rect 24861 4342 24907 4354
rect 24982 4676 25046 4688
rect 24982 4669 24997 4676
rect 25031 4669 25046 4676
rect 24982 4617 24988 4669
rect 25040 4617 25046 4669
rect 24982 4605 25046 4617
rect 24982 4553 24988 4605
rect 25040 4553 25046 4605
rect 24982 4541 25046 4553
rect 24982 4489 24988 4541
rect 25040 4489 25046 4541
rect 24982 4477 25046 4489
rect 24982 4425 24988 4477
rect 25040 4425 25046 4477
rect 24982 4413 25046 4425
rect 24982 4361 24988 4413
rect 25040 4361 25046 4413
rect 24982 4354 24997 4361
rect 25031 4354 25046 4361
rect 24982 4342 25046 4354
rect 25251 4676 25297 4902
rect 25381 5008 25427 5013
rect 25381 4974 25387 5008
rect 25421 4974 25427 5008
rect 25381 4936 25427 4974
rect 25381 4902 25387 4936
rect 25421 4902 25427 4936
rect 25381 4890 25427 4902
rect 25511 5008 25557 5013
rect 25511 4974 25517 5008
rect 25551 4974 25557 5008
rect 25511 4936 25557 4974
rect 25511 4902 25517 4936
rect 25551 4902 25557 4936
rect 25511 4890 25557 4902
rect 25641 5008 25687 5046
rect 25757 5089 25831 5113
rect 25757 5037 25768 5089
rect 25820 5037 25831 5089
rect 25757 5013 25831 5037
rect 25887 5089 25961 5113
rect 25887 5037 25898 5089
rect 25950 5037 25961 5089
rect 25887 5013 25961 5037
rect 26031 5080 26077 5118
rect 26161 5224 26207 5236
rect 26161 5190 26167 5224
rect 26201 5190 26207 5224
rect 26161 5152 26207 5190
rect 26161 5118 26167 5152
rect 26201 5118 26207 5152
rect 26161 5113 26207 5118
rect 26291 5224 26337 5236
rect 26291 5190 26297 5224
rect 26331 5190 26337 5224
rect 26291 5152 26337 5190
rect 26291 5118 26297 5152
rect 26331 5118 26337 5152
rect 26291 5113 26337 5118
rect 26421 5224 26467 5236
rect 26421 5190 26427 5224
rect 26461 5190 26467 5224
rect 26421 5152 26467 5190
rect 26421 5118 26427 5152
rect 26461 5118 26467 5152
rect 26031 5046 26037 5080
rect 26071 5046 26077 5080
rect 25641 4974 25647 5008
rect 25681 4974 25687 5008
rect 25641 4936 25687 4974
rect 25641 4902 25647 4936
rect 25681 4902 25687 4936
rect 25251 4642 25257 4676
rect 25291 4642 25297 4676
rect 25251 4604 25297 4642
rect 25251 4570 25257 4604
rect 25291 4570 25297 4604
rect 25251 4532 25297 4570
rect 25251 4498 25257 4532
rect 25291 4498 25297 4532
rect 25251 4460 25297 4498
rect 25251 4426 25257 4460
rect 25291 4426 25297 4460
rect 25251 4388 25297 4426
rect 25251 4354 25257 4388
rect 25291 4354 25297 4388
rect 25251 4342 25297 4354
rect 25372 4676 25436 4688
rect 25372 4669 25387 4676
rect 25421 4669 25436 4676
rect 25372 4617 25378 4669
rect 25430 4617 25436 4669
rect 25372 4605 25436 4617
rect 25372 4553 25378 4605
rect 25430 4553 25436 4605
rect 25372 4541 25436 4553
rect 25372 4489 25378 4541
rect 25430 4489 25436 4541
rect 25372 4477 25436 4489
rect 25372 4425 25378 4477
rect 25430 4425 25436 4477
rect 25372 4413 25436 4425
rect 25372 4361 25378 4413
rect 25430 4361 25436 4413
rect 25372 4354 25387 4361
rect 25421 4354 25436 4361
rect 25372 4342 25436 4354
rect 25641 4676 25687 4902
rect 25771 5008 25817 5013
rect 25771 4974 25777 5008
rect 25811 4974 25817 5008
rect 25771 4936 25817 4974
rect 25771 4902 25777 4936
rect 25811 4902 25817 4936
rect 25771 4890 25817 4902
rect 25901 5008 25947 5013
rect 25901 4974 25907 5008
rect 25941 4974 25947 5008
rect 25901 4936 25947 4974
rect 25901 4902 25907 4936
rect 25941 4902 25947 4936
rect 25901 4890 25947 4902
rect 26031 5008 26077 5046
rect 26147 5089 26221 5113
rect 26147 5037 26158 5089
rect 26210 5037 26221 5089
rect 26147 5013 26221 5037
rect 26277 5089 26351 5113
rect 26277 5037 26288 5089
rect 26340 5037 26351 5089
rect 26277 5013 26351 5037
rect 26421 5080 26467 5118
rect 26551 5224 26597 5236
rect 26551 5190 26557 5224
rect 26591 5190 26597 5224
rect 26551 5152 26597 5190
rect 26551 5118 26557 5152
rect 26591 5118 26597 5152
rect 26551 5113 26597 5118
rect 26681 5224 26727 5236
rect 26681 5190 26687 5224
rect 26721 5190 26727 5224
rect 26681 5152 26727 5190
rect 26681 5118 26687 5152
rect 26721 5118 26727 5152
rect 26681 5113 26727 5118
rect 26421 5046 26427 5080
rect 26461 5046 26467 5080
rect 26031 4974 26037 5008
rect 26071 4974 26077 5008
rect 26031 4936 26077 4974
rect 26031 4902 26037 4936
rect 26071 4902 26077 4936
rect 25641 4642 25647 4676
rect 25681 4642 25687 4676
rect 25641 4604 25687 4642
rect 25641 4570 25647 4604
rect 25681 4570 25687 4604
rect 25641 4532 25687 4570
rect 25641 4498 25647 4532
rect 25681 4498 25687 4532
rect 25641 4460 25687 4498
rect 25641 4426 25647 4460
rect 25681 4426 25687 4460
rect 25641 4388 25687 4426
rect 25641 4354 25647 4388
rect 25681 4354 25687 4388
rect 25641 4342 25687 4354
rect 25762 4676 25826 4688
rect 25762 4669 25777 4676
rect 25811 4669 25826 4676
rect 25762 4617 25768 4669
rect 25820 4617 25826 4669
rect 25762 4605 25826 4617
rect 25762 4553 25768 4605
rect 25820 4553 25826 4605
rect 25762 4541 25826 4553
rect 25762 4489 25768 4541
rect 25820 4489 25826 4541
rect 25762 4477 25826 4489
rect 25762 4425 25768 4477
rect 25820 4425 25826 4477
rect 25762 4413 25826 4425
rect 25762 4361 25768 4413
rect 25820 4361 25826 4413
rect 25762 4354 25777 4361
rect 25811 4354 25826 4361
rect 25762 4342 25826 4354
rect 26031 4676 26077 4902
rect 26161 5008 26207 5013
rect 26161 4974 26167 5008
rect 26201 4974 26207 5008
rect 26161 4936 26207 4974
rect 26161 4902 26167 4936
rect 26201 4902 26207 4936
rect 26161 4890 26207 4902
rect 26291 5008 26337 5013
rect 26291 4974 26297 5008
rect 26331 4974 26337 5008
rect 26291 4936 26337 4974
rect 26291 4902 26297 4936
rect 26331 4902 26337 4936
rect 26291 4890 26337 4902
rect 26421 5008 26467 5046
rect 26537 5089 26611 5113
rect 26537 5037 26548 5089
rect 26600 5037 26611 5089
rect 26537 5013 26611 5037
rect 26667 5089 26741 5113
rect 26667 5037 26678 5089
rect 26730 5037 26741 5089
rect 26667 5013 26741 5037
rect 26421 4974 26427 5008
rect 26461 4974 26467 5008
rect 26421 4936 26467 4974
rect 26421 4902 26427 4936
rect 26461 4902 26467 4936
rect 26031 4642 26037 4676
rect 26071 4642 26077 4676
rect 26031 4604 26077 4642
rect 26031 4570 26037 4604
rect 26071 4570 26077 4604
rect 26031 4532 26077 4570
rect 26031 4498 26037 4532
rect 26071 4498 26077 4532
rect 26031 4460 26077 4498
rect 26031 4426 26037 4460
rect 26071 4426 26077 4460
rect 26031 4388 26077 4426
rect 26031 4354 26037 4388
rect 26071 4354 26077 4388
rect 26031 4342 26077 4354
rect 26152 4676 26216 4688
rect 26152 4669 26167 4676
rect 26201 4669 26216 4676
rect 26152 4617 26158 4669
rect 26210 4617 26216 4669
rect 26152 4605 26216 4617
rect 26152 4553 26158 4605
rect 26210 4553 26216 4605
rect 26152 4541 26216 4553
rect 26152 4489 26158 4541
rect 26210 4489 26216 4541
rect 26152 4477 26216 4489
rect 26152 4425 26158 4477
rect 26210 4425 26216 4477
rect 26152 4413 26216 4425
rect 26152 4361 26158 4413
rect 26210 4361 26216 4413
rect 26152 4354 26167 4361
rect 26201 4354 26216 4361
rect 26152 4342 26216 4354
rect 26421 4676 26467 4902
rect 26551 5008 26597 5013
rect 26551 4974 26557 5008
rect 26591 4974 26597 5008
rect 26551 4936 26597 4974
rect 26551 4902 26557 4936
rect 26591 4902 26597 4936
rect 26551 4890 26597 4902
rect 26681 5008 26727 5013
rect 26681 4974 26687 5008
rect 26721 4974 26727 5008
rect 26681 4936 26727 4974
rect 26681 4902 26687 4936
rect 26721 4902 26727 4936
rect 26681 4890 26727 4902
rect 26876 4924 27116 4927
rect 26876 4915 26909 4924
rect 26876 4881 26907 4915
rect 26876 4872 26909 4881
rect 26961 4872 26973 4924
rect 27025 4872 27037 4924
rect 27089 4872 27116 4924
rect 26876 4869 27116 4872
rect 26790 4781 26796 4833
rect 26848 4827 26854 4833
rect 26967 4827 27127 4834
rect 26848 4824 27127 4827
rect 26848 4790 26994 4824
rect 27028 4790 27066 4824
rect 27100 4790 27127 4824
rect 26848 4787 27127 4790
rect 26848 4781 26854 4787
rect 26967 4780 27127 4787
rect 26421 4642 26427 4676
rect 26461 4642 26467 4676
rect 26421 4604 26467 4642
rect 26421 4570 26427 4604
rect 26461 4570 26467 4604
rect 26421 4532 26467 4570
rect 26421 4498 26427 4532
rect 26461 4498 26467 4532
rect 26421 4460 26467 4498
rect 26421 4426 26427 4460
rect 26461 4426 26467 4460
rect 26421 4388 26467 4426
rect 26421 4354 26427 4388
rect 26461 4354 26467 4388
rect 26421 4342 26467 4354
rect 26542 4676 26606 4688
rect 26542 4669 26557 4676
rect 26591 4669 26606 4676
rect 26542 4617 26548 4669
rect 26600 4617 26606 4669
rect 26542 4605 26606 4617
rect 26542 4553 26548 4605
rect 26600 4553 26606 4605
rect 26542 4541 26606 4553
rect 26542 4489 26548 4541
rect 26600 4489 26606 4541
rect 26542 4477 26606 4489
rect 26542 4425 26548 4477
rect 26600 4425 26606 4477
rect 26542 4413 26606 4425
rect 26542 4361 26548 4413
rect 26600 4361 26606 4413
rect 26795 4676 26841 4688
rect 26885 4685 26931 4688
rect 26795 4642 26801 4676
rect 26835 4642 26841 4676
rect 26795 4604 26841 4642
rect 26876 4633 26882 4685
rect 26934 4633 26940 4685
rect 26975 4676 27021 4688
rect 27065 4685 27111 4688
rect 26975 4642 26981 4676
rect 27015 4642 27021 4676
rect 26795 4570 26801 4604
rect 26835 4570 26841 4604
rect 26795 4532 26841 4570
rect 26795 4498 26801 4532
rect 26835 4498 26841 4532
rect 26795 4460 26841 4498
rect 26795 4426 26801 4460
rect 26835 4426 26841 4460
rect 26795 4397 26841 4426
rect 26885 4604 26931 4633
rect 26885 4570 26891 4604
rect 26925 4570 26931 4604
rect 26885 4532 26931 4570
rect 26885 4498 26891 4532
rect 26925 4498 26931 4532
rect 26885 4460 26931 4498
rect 26885 4426 26891 4460
rect 26925 4426 26931 4460
rect 26542 4354 26557 4361
rect 26591 4354 26606 4361
rect 26542 4342 26606 4354
rect 26786 4345 26792 4397
rect 26844 4345 26850 4397
rect 26885 4388 26931 4426
rect 26975 4604 27021 4642
rect 27056 4633 27062 4685
rect 27114 4633 27120 4685
rect 27155 4676 27201 4688
rect 27155 4642 27161 4676
rect 27195 4642 27201 4676
rect 26975 4570 26981 4604
rect 27015 4570 27021 4604
rect 26975 4532 27021 4570
rect 26975 4498 26981 4532
rect 27015 4498 27021 4532
rect 26975 4460 27021 4498
rect 26975 4426 26981 4460
rect 27015 4426 27021 4460
rect 26975 4392 27021 4426
rect 27065 4604 27111 4633
rect 27065 4570 27071 4604
rect 27105 4570 27111 4604
rect 27065 4532 27111 4570
rect 27065 4498 27071 4532
rect 27105 4498 27111 4532
rect 27065 4460 27111 4498
rect 27065 4426 27071 4460
rect 27105 4426 27111 4460
rect 26885 4354 26891 4388
rect 26925 4354 26931 4388
rect 26795 4342 26841 4345
rect 26885 4342 26931 4354
rect 26965 4391 27031 4392
rect 15553 4338 15619 4339
rect 26965 4339 26972 4391
rect 27024 4339 27031 4391
rect 27065 4388 27111 4426
rect 27155 4604 27201 4642
rect 27155 4570 27161 4604
rect 27195 4570 27201 4604
rect 27155 4532 27201 4570
rect 27155 4498 27161 4532
rect 27195 4498 27201 4532
rect 27155 4460 27201 4498
rect 27155 4426 27161 4460
rect 27195 4426 27201 4460
rect 27155 4392 27201 4426
rect 27065 4354 27071 4388
rect 27105 4354 27111 4388
rect 27065 4342 27111 4354
rect 27145 4391 27211 4392
rect 26965 4338 27031 4339
rect 27145 4339 27152 4391
rect 27204 4339 27211 4391
rect 27145 4338 27211 4339
rect 15797 4296 15957 4302
rect 27389 4296 27549 4302
rect 15373 4295 15957 4296
rect 15373 4243 15380 4295
rect 15432 4243 15560 4295
rect 15612 4243 15819 4295
rect 15871 4243 15883 4295
rect 15935 4243 15957 4295
rect 15373 4242 15957 4243
rect 26965 4295 27549 4296
rect 26965 4243 26972 4295
rect 27024 4243 27152 4295
rect 27204 4243 27411 4295
rect 27463 4243 27475 4295
rect 27527 4243 27549 4295
rect 26965 4242 27549 4243
rect 15797 4236 15957 4242
rect 27389 4236 27549 4242
rect 12891 4117 13294 4123
rect 12891 4065 12897 4117
rect 12949 4108 13294 4117
rect 12949 4074 13244 4108
rect 13278 4074 13294 4108
rect 12949 4065 13294 4074
rect 12891 4059 13294 4065
rect 13390 4117 13684 4123
rect 13390 4065 13396 4117
rect 13448 4108 13684 4117
rect 13448 4074 13634 4108
rect 13668 4074 13684 4108
rect 13448 4065 13684 4074
rect 13390 4059 13684 4065
rect 13780 4117 14074 4123
rect 13780 4065 13786 4117
rect 13838 4108 14074 4117
rect 13838 4074 14024 4108
rect 14058 4074 14074 4108
rect 13838 4065 14074 4074
rect 13780 4059 14074 4065
rect 14170 4117 14464 4123
rect 14170 4065 14176 4117
rect 14228 4108 14464 4117
rect 14228 4074 14414 4108
rect 14448 4074 14464 4108
rect 14228 4065 14464 4074
rect 14170 4059 14464 4065
rect 14560 4117 14854 4123
rect 14560 4065 14566 4117
rect 14618 4108 14854 4117
rect 14618 4074 14804 4108
rect 14838 4074 14854 4108
rect 14618 4065 14854 4074
rect 14560 4059 14854 4065
rect 14950 4117 15729 4123
rect 14950 4065 14956 4117
rect 15008 4108 15671 4117
rect 15008 4074 15249 4108
rect 15283 4074 15671 4108
rect 15008 4065 15671 4074
rect 15723 4065 15729 4117
rect 14950 4059 15729 4065
rect 24483 4117 24886 4123
rect 24483 4065 24489 4117
rect 24541 4108 24886 4117
rect 24541 4074 24836 4108
rect 24870 4074 24886 4108
rect 24541 4065 24886 4074
rect 24483 4059 24886 4065
rect 24982 4117 25276 4123
rect 24982 4065 24988 4117
rect 25040 4108 25276 4117
rect 25040 4074 25226 4108
rect 25260 4074 25276 4108
rect 25040 4065 25276 4074
rect 24982 4059 25276 4065
rect 25372 4117 25666 4123
rect 25372 4065 25378 4117
rect 25430 4108 25666 4117
rect 25430 4074 25616 4108
rect 25650 4074 25666 4108
rect 25430 4065 25666 4074
rect 25372 4059 25666 4065
rect 25762 4117 26056 4123
rect 25762 4065 25768 4117
rect 25820 4108 26056 4117
rect 25820 4074 26006 4108
rect 26040 4074 26056 4108
rect 25820 4065 26056 4074
rect 25762 4059 26056 4065
rect 26152 4117 26446 4123
rect 26152 4065 26158 4117
rect 26210 4108 26446 4117
rect 26210 4074 26396 4108
rect 26430 4074 26446 4108
rect 26210 4065 26446 4074
rect 26152 4059 26446 4065
rect 26542 4117 27321 4123
rect 26542 4065 26548 4117
rect 26600 4108 27263 4117
rect 26600 4074 26841 4108
rect 26875 4074 27263 4108
rect 26600 4065 27263 4074
rect 27315 4065 27321 4117
rect 26542 4059 27321 4065
rect 12590 3960 15729 3961
rect 12590 3908 12596 3960
rect 12648 3951 15729 3960
rect 12648 3917 13860 3951
rect 13894 3917 14640 3951
rect 14674 3917 15729 3951
rect 12648 3908 15729 3917
rect 12590 3907 15729 3908
rect 24182 3960 27321 3961
rect 24182 3908 24188 3960
rect 24240 3951 27321 3960
rect 24240 3917 25452 3951
rect 25486 3917 26232 3951
rect 26266 3917 27321 3951
rect 24240 3908 27321 3917
rect 24182 3907 27321 3908
rect 13269 3820 13315 3832
rect 13269 3786 13275 3820
rect 13309 3786 13315 3820
rect 13269 3748 13315 3786
rect 13269 3714 13275 3748
rect 13309 3714 13315 3748
rect 13000 3477 13064 3484
rect 13000 3425 13006 3477
rect 13058 3425 13064 3477
rect 13139 3472 13185 3484
rect 13139 3469 13145 3472
rect 13000 3413 13064 3425
rect 12585 3398 12659 3405
rect 12585 3346 12596 3398
rect 12648 3346 12659 3398
rect 13000 3361 13006 3413
rect 13058 3361 13064 3413
rect 13125 3445 13145 3469
rect 13179 3469 13185 3472
rect 13269 3472 13315 3714
rect 13390 3825 13454 3832
rect 13390 3773 13396 3825
rect 13448 3773 13454 3825
rect 13390 3761 13454 3773
rect 13390 3709 13396 3761
rect 13448 3709 13454 3761
rect 13390 3702 13454 3709
rect 13520 3825 13584 3832
rect 13520 3773 13526 3825
rect 13578 3773 13584 3825
rect 13520 3761 13584 3773
rect 13520 3709 13526 3761
rect 13578 3709 13584 3761
rect 13520 3702 13584 3709
rect 13659 3820 13705 3832
rect 13659 3786 13665 3820
rect 13699 3786 13705 3820
rect 13659 3748 13705 3786
rect 13659 3714 13665 3748
rect 13699 3714 13705 3748
rect 13179 3445 13199 3469
rect 13125 3393 13136 3445
rect 13188 3393 13199 3445
rect 13125 3369 13145 3393
rect 13000 3354 13064 3361
rect 13139 3366 13145 3369
rect 13179 3369 13199 3393
rect 13269 3438 13275 3472
rect 13309 3438 13315 3472
rect 13399 3472 13445 3484
rect 13399 3469 13405 3472
rect 13269 3400 13315 3438
rect 13179 3366 13185 3369
rect 13139 3354 13185 3366
rect 13269 3366 13275 3400
rect 13309 3366 13315 3400
rect 13385 3445 13405 3469
rect 13439 3469 13445 3472
rect 13529 3472 13575 3484
rect 13529 3469 13535 3472
rect 13439 3445 13459 3469
rect 13385 3393 13396 3445
rect 13448 3393 13459 3445
rect 13385 3369 13405 3393
rect 13269 3354 13315 3366
rect 13399 3366 13405 3369
rect 13439 3369 13459 3393
rect 13515 3445 13535 3469
rect 13569 3469 13575 3472
rect 13659 3472 13705 3714
rect 13780 3825 13844 3832
rect 13780 3773 13786 3825
rect 13838 3773 13844 3825
rect 13780 3761 13844 3773
rect 13780 3709 13786 3761
rect 13838 3709 13844 3761
rect 13780 3702 13844 3709
rect 13910 3825 13974 3832
rect 13910 3773 13916 3825
rect 13968 3773 13974 3825
rect 13910 3761 13974 3773
rect 13910 3709 13916 3761
rect 13968 3709 13974 3761
rect 13910 3702 13974 3709
rect 14049 3820 14095 3832
rect 14049 3786 14055 3820
rect 14089 3786 14095 3820
rect 14049 3748 14095 3786
rect 14049 3714 14055 3748
rect 14089 3714 14095 3748
rect 13569 3445 13589 3469
rect 13515 3393 13526 3445
rect 13578 3393 13589 3445
rect 13515 3369 13535 3393
rect 13439 3366 13445 3369
rect 13399 3354 13445 3366
rect 13529 3366 13535 3369
rect 13569 3369 13589 3393
rect 13659 3438 13665 3472
rect 13699 3438 13705 3472
rect 13789 3472 13835 3484
rect 13789 3469 13795 3472
rect 13659 3400 13705 3438
rect 13569 3366 13575 3369
rect 13529 3354 13575 3366
rect 13659 3366 13665 3400
rect 13699 3366 13705 3400
rect 13775 3445 13795 3469
rect 13829 3469 13835 3472
rect 13919 3472 13965 3484
rect 13919 3469 13925 3472
rect 13829 3445 13849 3469
rect 13775 3393 13786 3445
rect 13838 3393 13849 3445
rect 13775 3369 13795 3393
rect 13659 3354 13705 3366
rect 13789 3366 13795 3369
rect 13829 3369 13849 3393
rect 13905 3445 13925 3469
rect 13959 3469 13965 3472
rect 14049 3472 14095 3714
rect 14170 3825 14234 3832
rect 14170 3773 14176 3825
rect 14228 3773 14234 3825
rect 14170 3761 14234 3773
rect 14170 3709 14176 3761
rect 14228 3709 14234 3761
rect 14170 3702 14234 3709
rect 14300 3825 14364 3832
rect 14300 3773 14306 3825
rect 14358 3773 14364 3825
rect 14300 3761 14364 3773
rect 14300 3709 14306 3761
rect 14358 3709 14364 3761
rect 14300 3702 14364 3709
rect 14439 3820 14485 3832
rect 14439 3786 14445 3820
rect 14479 3786 14485 3820
rect 14439 3748 14485 3786
rect 14439 3714 14445 3748
rect 14479 3714 14485 3748
rect 13959 3445 13979 3469
rect 13905 3393 13916 3445
rect 13968 3393 13979 3445
rect 13905 3369 13925 3393
rect 13829 3366 13835 3369
rect 13789 3354 13835 3366
rect 13919 3366 13925 3369
rect 13959 3369 13979 3393
rect 14049 3438 14055 3472
rect 14089 3438 14095 3472
rect 14179 3472 14225 3484
rect 14179 3469 14185 3472
rect 14049 3400 14095 3438
rect 13959 3366 13965 3369
rect 13919 3354 13965 3366
rect 14049 3366 14055 3400
rect 14089 3366 14095 3400
rect 14165 3445 14185 3469
rect 14219 3469 14225 3472
rect 14309 3472 14355 3484
rect 14309 3469 14315 3472
rect 14219 3445 14239 3469
rect 14165 3393 14176 3445
rect 14228 3393 14239 3445
rect 14165 3369 14185 3393
rect 14049 3354 14095 3366
rect 14179 3366 14185 3369
rect 14219 3369 14239 3393
rect 14295 3445 14315 3469
rect 14349 3469 14355 3472
rect 14439 3472 14485 3714
rect 14560 3825 14624 3832
rect 14560 3773 14566 3825
rect 14618 3773 14624 3825
rect 14560 3761 14624 3773
rect 14560 3709 14566 3761
rect 14618 3709 14624 3761
rect 14560 3702 14624 3709
rect 14690 3825 14754 3832
rect 14690 3773 14696 3825
rect 14748 3773 14754 3825
rect 14690 3761 14754 3773
rect 14690 3709 14696 3761
rect 14748 3709 14754 3761
rect 14690 3702 14754 3709
rect 14829 3820 14875 3832
rect 14829 3786 14835 3820
rect 14869 3786 14875 3820
rect 14829 3748 14875 3786
rect 14829 3714 14835 3748
rect 14869 3714 14875 3748
rect 14349 3445 14369 3469
rect 14295 3393 14306 3445
rect 14358 3393 14369 3445
rect 14295 3369 14315 3393
rect 14219 3366 14225 3369
rect 14179 3354 14225 3366
rect 14309 3366 14315 3369
rect 14349 3369 14369 3393
rect 14439 3438 14445 3472
rect 14479 3438 14485 3472
rect 14569 3472 14615 3484
rect 14569 3469 14575 3472
rect 14439 3400 14485 3438
rect 14349 3366 14355 3369
rect 14309 3354 14355 3366
rect 14439 3366 14445 3400
rect 14479 3366 14485 3400
rect 14555 3445 14575 3469
rect 14609 3469 14615 3472
rect 14699 3472 14745 3484
rect 14699 3469 14705 3472
rect 14609 3445 14629 3469
rect 14555 3393 14566 3445
rect 14618 3393 14629 3445
rect 14555 3369 14575 3393
rect 14439 3354 14485 3366
rect 14569 3366 14575 3369
rect 14609 3369 14629 3393
rect 14685 3445 14705 3469
rect 14739 3469 14745 3472
rect 14829 3472 14875 3714
rect 14950 3825 15014 3832
rect 14950 3773 14956 3825
rect 15008 3773 15014 3825
rect 14950 3761 15014 3773
rect 14950 3709 14956 3761
rect 15008 3709 15014 3761
rect 14950 3702 15014 3709
rect 15080 3825 15144 3832
rect 15203 3829 15249 3832
rect 15080 3773 15086 3825
rect 15138 3773 15144 3825
rect 15194 3777 15200 3829
rect 15252 3777 15258 3829
rect 15293 3820 15339 3832
rect 15383 3829 15429 3832
rect 15293 3786 15299 3820
rect 15333 3786 15339 3820
rect 15080 3761 15144 3773
rect 15080 3709 15086 3761
rect 15138 3709 15144 3761
rect 15080 3702 15144 3709
rect 15203 3748 15249 3777
rect 15293 3757 15339 3786
rect 15374 3777 15380 3829
rect 15432 3777 15438 3829
rect 15473 3820 15519 3832
rect 15563 3829 15609 3832
rect 15473 3786 15479 3820
rect 15513 3786 15519 3820
rect 15203 3714 15209 3748
rect 15243 3714 15249 3748
rect 15203 3702 15249 3714
rect 15284 3705 15290 3757
rect 15342 3705 15348 3757
rect 15383 3748 15429 3777
rect 15473 3757 15519 3786
rect 15554 3777 15560 3829
rect 15612 3777 15618 3829
rect 24861 3820 24907 3832
rect 24861 3786 24867 3820
rect 24901 3786 24907 3820
rect 15383 3714 15389 3748
rect 15423 3714 15429 3748
rect 15293 3702 15339 3705
rect 15383 3702 15429 3714
rect 15464 3705 15470 3757
rect 15522 3705 15528 3757
rect 15563 3748 15609 3777
rect 15563 3714 15569 3748
rect 15603 3714 15609 3748
rect 15473 3702 15519 3705
rect 15563 3702 15609 3714
rect 24861 3748 24907 3786
rect 24861 3714 24867 3748
rect 24901 3714 24907 3748
rect 15287 3588 15527 3591
rect 15287 3536 15316 3588
rect 15368 3536 15380 3588
rect 15432 3536 15444 3588
rect 15496 3536 15527 3588
rect 15287 3533 15527 3536
rect 14739 3445 14759 3469
rect 14685 3393 14696 3445
rect 14748 3393 14759 3445
rect 14685 3369 14705 3393
rect 14609 3366 14615 3369
rect 14569 3354 14615 3366
rect 14699 3366 14705 3369
rect 14739 3369 14759 3393
rect 14829 3438 14835 3472
rect 14869 3438 14875 3472
rect 14959 3472 15005 3484
rect 14959 3469 14965 3472
rect 14829 3400 14875 3438
rect 14739 3366 14745 3369
rect 14699 3354 14745 3366
rect 14829 3366 14835 3400
rect 14869 3366 14875 3400
rect 14945 3445 14965 3469
rect 14999 3469 15005 3472
rect 15089 3472 15135 3484
rect 15089 3469 15095 3472
rect 14999 3445 15019 3469
rect 14945 3393 14956 3445
rect 15008 3393 15019 3445
rect 14945 3369 14965 3393
rect 14829 3354 14875 3366
rect 14959 3366 14965 3369
rect 14999 3369 15019 3393
rect 15075 3445 15095 3469
rect 15129 3469 15135 3472
rect 24592 3477 24656 3484
rect 15129 3445 15149 3469
rect 15075 3393 15086 3445
rect 15138 3393 15149 3445
rect 24592 3425 24598 3477
rect 24650 3425 24656 3477
rect 24731 3472 24777 3484
rect 24731 3469 24737 3472
rect 24592 3413 24656 3425
rect 15075 3369 15095 3393
rect 14999 3366 15005 3369
rect 14959 3354 15005 3366
rect 15089 3366 15095 3369
rect 15129 3369 15149 3393
rect 24177 3398 24251 3405
rect 15129 3366 15135 3369
rect 15089 3354 15135 3366
rect 12585 3339 12659 3346
rect 24177 3346 24188 3398
rect 24240 3346 24251 3398
rect 24592 3361 24598 3413
rect 24650 3361 24656 3413
rect 24717 3445 24737 3469
rect 24771 3469 24777 3472
rect 24861 3472 24907 3714
rect 24982 3825 25046 3832
rect 24982 3773 24988 3825
rect 25040 3773 25046 3825
rect 24982 3761 25046 3773
rect 24982 3709 24988 3761
rect 25040 3709 25046 3761
rect 24982 3702 25046 3709
rect 25112 3825 25176 3832
rect 25112 3773 25118 3825
rect 25170 3773 25176 3825
rect 25112 3761 25176 3773
rect 25112 3709 25118 3761
rect 25170 3709 25176 3761
rect 25112 3702 25176 3709
rect 25251 3820 25297 3832
rect 25251 3786 25257 3820
rect 25291 3786 25297 3820
rect 25251 3748 25297 3786
rect 25251 3714 25257 3748
rect 25291 3714 25297 3748
rect 24771 3445 24791 3469
rect 24717 3393 24728 3445
rect 24780 3393 24791 3445
rect 24717 3369 24737 3393
rect 24592 3354 24656 3361
rect 24731 3366 24737 3369
rect 24771 3369 24791 3393
rect 24861 3438 24867 3472
rect 24901 3438 24907 3472
rect 24991 3472 25037 3484
rect 24991 3469 24997 3472
rect 24861 3400 24907 3438
rect 24771 3366 24777 3369
rect 24731 3354 24777 3366
rect 24861 3366 24867 3400
rect 24901 3366 24907 3400
rect 24977 3445 24997 3469
rect 25031 3469 25037 3472
rect 25121 3472 25167 3484
rect 25121 3469 25127 3472
rect 25031 3445 25051 3469
rect 24977 3393 24988 3445
rect 25040 3393 25051 3445
rect 24977 3369 24997 3393
rect 24861 3354 24907 3366
rect 24991 3366 24997 3369
rect 25031 3369 25051 3393
rect 25107 3445 25127 3469
rect 25161 3469 25167 3472
rect 25251 3472 25297 3714
rect 25372 3825 25436 3832
rect 25372 3773 25378 3825
rect 25430 3773 25436 3825
rect 25372 3761 25436 3773
rect 25372 3709 25378 3761
rect 25430 3709 25436 3761
rect 25372 3702 25436 3709
rect 25502 3825 25566 3832
rect 25502 3773 25508 3825
rect 25560 3773 25566 3825
rect 25502 3761 25566 3773
rect 25502 3709 25508 3761
rect 25560 3709 25566 3761
rect 25502 3702 25566 3709
rect 25641 3820 25687 3832
rect 25641 3786 25647 3820
rect 25681 3786 25687 3820
rect 25641 3748 25687 3786
rect 25641 3714 25647 3748
rect 25681 3714 25687 3748
rect 25161 3445 25181 3469
rect 25107 3393 25118 3445
rect 25170 3393 25181 3445
rect 25107 3369 25127 3393
rect 25031 3366 25037 3369
rect 24991 3354 25037 3366
rect 25121 3366 25127 3369
rect 25161 3369 25181 3393
rect 25251 3438 25257 3472
rect 25291 3438 25297 3472
rect 25381 3472 25427 3484
rect 25381 3469 25387 3472
rect 25251 3400 25297 3438
rect 25161 3366 25167 3369
rect 25121 3354 25167 3366
rect 25251 3366 25257 3400
rect 25291 3366 25297 3400
rect 25367 3445 25387 3469
rect 25421 3469 25427 3472
rect 25511 3472 25557 3484
rect 25511 3469 25517 3472
rect 25421 3445 25441 3469
rect 25367 3393 25378 3445
rect 25430 3393 25441 3445
rect 25367 3369 25387 3393
rect 25251 3354 25297 3366
rect 25381 3366 25387 3369
rect 25421 3369 25441 3393
rect 25497 3445 25517 3469
rect 25551 3469 25557 3472
rect 25641 3472 25687 3714
rect 25762 3825 25826 3832
rect 25762 3773 25768 3825
rect 25820 3773 25826 3825
rect 25762 3761 25826 3773
rect 25762 3709 25768 3761
rect 25820 3709 25826 3761
rect 25762 3702 25826 3709
rect 25892 3825 25956 3832
rect 25892 3773 25898 3825
rect 25950 3773 25956 3825
rect 25892 3761 25956 3773
rect 25892 3709 25898 3761
rect 25950 3709 25956 3761
rect 25892 3702 25956 3709
rect 26031 3820 26077 3832
rect 26031 3786 26037 3820
rect 26071 3786 26077 3820
rect 26031 3748 26077 3786
rect 26031 3714 26037 3748
rect 26071 3714 26077 3748
rect 25551 3445 25571 3469
rect 25497 3393 25508 3445
rect 25560 3393 25571 3445
rect 25497 3369 25517 3393
rect 25421 3366 25427 3369
rect 25381 3354 25427 3366
rect 25511 3366 25517 3369
rect 25551 3369 25571 3393
rect 25641 3438 25647 3472
rect 25681 3438 25687 3472
rect 25771 3472 25817 3484
rect 25771 3469 25777 3472
rect 25641 3400 25687 3438
rect 25551 3366 25557 3369
rect 25511 3354 25557 3366
rect 25641 3366 25647 3400
rect 25681 3366 25687 3400
rect 25757 3445 25777 3469
rect 25811 3469 25817 3472
rect 25901 3472 25947 3484
rect 25901 3469 25907 3472
rect 25811 3445 25831 3469
rect 25757 3393 25768 3445
rect 25820 3393 25831 3445
rect 25757 3369 25777 3393
rect 25641 3354 25687 3366
rect 25771 3366 25777 3369
rect 25811 3369 25831 3393
rect 25887 3445 25907 3469
rect 25941 3469 25947 3472
rect 26031 3472 26077 3714
rect 26152 3825 26216 3832
rect 26152 3773 26158 3825
rect 26210 3773 26216 3825
rect 26152 3761 26216 3773
rect 26152 3709 26158 3761
rect 26210 3709 26216 3761
rect 26152 3702 26216 3709
rect 26282 3825 26346 3832
rect 26282 3773 26288 3825
rect 26340 3773 26346 3825
rect 26282 3761 26346 3773
rect 26282 3709 26288 3761
rect 26340 3709 26346 3761
rect 26282 3702 26346 3709
rect 26421 3820 26467 3832
rect 26421 3786 26427 3820
rect 26461 3786 26467 3820
rect 26421 3748 26467 3786
rect 26421 3714 26427 3748
rect 26461 3714 26467 3748
rect 25941 3445 25961 3469
rect 25887 3393 25898 3445
rect 25950 3393 25961 3445
rect 25887 3369 25907 3393
rect 25811 3366 25817 3369
rect 25771 3354 25817 3366
rect 25901 3366 25907 3369
rect 25941 3369 25961 3393
rect 26031 3438 26037 3472
rect 26071 3438 26077 3472
rect 26161 3472 26207 3484
rect 26161 3469 26167 3472
rect 26031 3400 26077 3438
rect 25941 3366 25947 3369
rect 25901 3354 25947 3366
rect 26031 3366 26037 3400
rect 26071 3366 26077 3400
rect 26147 3445 26167 3469
rect 26201 3469 26207 3472
rect 26291 3472 26337 3484
rect 26291 3469 26297 3472
rect 26201 3445 26221 3469
rect 26147 3393 26158 3445
rect 26210 3393 26221 3445
rect 26147 3369 26167 3393
rect 26031 3354 26077 3366
rect 26161 3366 26167 3369
rect 26201 3369 26221 3393
rect 26277 3445 26297 3469
rect 26331 3469 26337 3472
rect 26421 3472 26467 3714
rect 26542 3825 26606 3832
rect 26542 3773 26548 3825
rect 26600 3773 26606 3825
rect 26542 3761 26606 3773
rect 26542 3709 26548 3761
rect 26600 3709 26606 3761
rect 26542 3702 26606 3709
rect 26672 3825 26736 3832
rect 26795 3829 26841 3832
rect 26672 3773 26678 3825
rect 26730 3773 26736 3825
rect 26786 3777 26792 3829
rect 26844 3777 26850 3829
rect 26885 3820 26931 3832
rect 26975 3829 27021 3832
rect 26885 3786 26891 3820
rect 26925 3786 26931 3820
rect 26672 3761 26736 3773
rect 26672 3709 26678 3761
rect 26730 3709 26736 3761
rect 26672 3702 26736 3709
rect 26795 3748 26841 3777
rect 26885 3757 26931 3786
rect 26966 3777 26972 3829
rect 27024 3777 27030 3829
rect 27065 3820 27111 3832
rect 27155 3829 27201 3832
rect 27065 3786 27071 3820
rect 27105 3786 27111 3820
rect 26795 3714 26801 3748
rect 26835 3714 26841 3748
rect 26795 3702 26841 3714
rect 26876 3705 26882 3757
rect 26934 3705 26940 3757
rect 26975 3748 27021 3777
rect 27065 3757 27111 3786
rect 27146 3777 27152 3829
rect 27204 3777 27210 3829
rect 26975 3714 26981 3748
rect 27015 3714 27021 3748
rect 26885 3702 26931 3705
rect 26975 3702 27021 3714
rect 27056 3705 27062 3757
rect 27114 3705 27120 3757
rect 27155 3748 27201 3777
rect 27155 3714 27161 3748
rect 27195 3714 27201 3748
rect 27065 3702 27111 3705
rect 27155 3702 27201 3714
rect 26879 3588 27119 3591
rect 26879 3536 26908 3588
rect 26960 3536 26972 3588
rect 27024 3536 27036 3588
rect 27088 3536 27119 3588
rect 26879 3533 27119 3536
rect 26331 3445 26351 3469
rect 26277 3393 26288 3445
rect 26340 3393 26351 3445
rect 26277 3369 26297 3393
rect 26201 3366 26207 3369
rect 26161 3354 26207 3366
rect 26291 3366 26297 3369
rect 26331 3369 26351 3393
rect 26421 3438 26427 3472
rect 26461 3438 26467 3472
rect 26551 3472 26597 3484
rect 26551 3469 26557 3472
rect 26421 3400 26467 3438
rect 26331 3366 26337 3369
rect 26291 3354 26337 3366
rect 26421 3366 26427 3400
rect 26461 3366 26467 3400
rect 26537 3445 26557 3469
rect 26591 3469 26597 3472
rect 26681 3472 26727 3484
rect 26681 3469 26687 3472
rect 26591 3445 26611 3469
rect 26537 3393 26548 3445
rect 26600 3393 26611 3445
rect 26537 3369 26557 3393
rect 26421 3354 26467 3366
rect 26551 3366 26557 3369
rect 26591 3369 26611 3393
rect 26667 3445 26687 3469
rect 26721 3469 26727 3472
rect 26721 3445 26741 3469
rect 26667 3393 26678 3445
rect 26730 3393 26741 3445
rect 26667 3369 26687 3393
rect 26591 3366 26597 3369
rect 26551 3354 26597 3366
rect 26681 3366 26687 3369
rect 26721 3369 26741 3393
rect 26721 3366 26727 3369
rect 26681 3354 26727 3366
rect 24177 3339 24251 3346
rect 12677 3272 12751 3279
rect 12677 3220 12688 3272
rect 12740 3220 12751 3272
rect 12677 3213 12751 3220
rect 12992 3272 13066 3279
rect 12992 3220 13003 3272
rect 13055 3220 13066 3272
rect 13320 3272 13394 3279
rect 12992 3213 13066 3220
rect 13190 3263 13264 3269
rect 13190 3229 13210 3263
rect 13244 3229 13264 3263
rect 13190 3153 13264 3229
rect 13320 3220 13331 3272
rect 13383 3220 13394 3272
rect 13710 3272 13784 3279
rect 13320 3213 13394 3220
rect 13450 3263 13524 3269
rect 13450 3229 13470 3263
rect 13504 3229 13524 3263
rect 13450 3153 13524 3229
rect 13580 3263 13654 3269
rect 13580 3229 13600 3263
rect 13634 3229 13654 3263
rect 13580 3153 13654 3229
rect 13710 3220 13721 3272
rect 13773 3220 13784 3272
rect 14100 3272 14174 3279
rect 13710 3213 13784 3220
rect 13840 3263 13914 3269
rect 13840 3229 13860 3263
rect 13894 3229 13914 3263
rect 13840 3153 13914 3229
rect 13970 3263 14044 3269
rect 13970 3229 13990 3263
rect 14024 3229 14044 3263
rect 13970 3153 14044 3229
rect 14100 3220 14111 3272
rect 14163 3220 14174 3272
rect 14490 3272 14564 3279
rect 14100 3213 14174 3220
rect 14230 3263 14304 3269
rect 14230 3229 14250 3263
rect 14284 3229 14304 3263
rect 14230 3153 14304 3229
rect 14360 3263 14434 3269
rect 14360 3229 14380 3263
rect 14414 3229 14434 3263
rect 14360 3153 14434 3229
rect 14490 3220 14501 3272
rect 14553 3220 14564 3272
rect 14880 3272 14954 3279
rect 14490 3213 14564 3220
rect 14620 3263 14694 3269
rect 14620 3229 14640 3263
rect 14674 3229 14694 3263
rect 14620 3153 14694 3229
rect 14750 3263 14824 3269
rect 14750 3229 14770 3263
rect 14804 3229 14824 3263
rect 14750 3153 14824 3229
rect 14880 3220 14891 3272
rect 14943 3220 14954 3272
rect 24269 3272 24343 3279
rect 14880 3213 14954 3220
rect 15010 3263 15084 3269
rect 15010 3229 15030 3263
rect 15064 3229 15084 3263
rect 15010 3153 15084 3229
rect 24269 3220 24280 3272
rect 24332 3220 24343 3272
rect 24269 3213 24343 3220
rect 24584 3272 24658 3279
rect 24584 3220 24595 3272
rect 24647 3220 24658 3272
rect 24912 3272 24986 3279
rect 24584 3213 24658 3220
rect 24782 3263 24856 3269
rect 24782 3229 24802 3263
rect 24836 3229 24856 3263
rect 24782 3153 24856 3229
rect 24912 3220 24923 3272
rect 24975 3220 24986 3272
rect 25302 3272 25376 3279
rect 24912 3213 24986 3220
rect 25042 3263 25116 3269
rect 25042 3229 25062 3263
rect 25096 3229 25116 3263
rect 25042 3153 25116 3229
rect 25172 3263 25246 3269
rect 25172 3229 25192 3263
rect 25226 3229 25246 3263
rect 25172 3153 25246 3229
rect 25302 3220 25313 3272
rect 25365 3220 25376 3272
rect 25692 3272 25766 3279
rect 25302 3213 25376 3220
rect 25432 3263 25506 3269
rect 25432 3229 25452 3263
rect 25486 3229 25506 3263
rect 25432 3153 25506 3229
rect 25562 3263 25636 3269
rect 25562 3229 25582 3263
rect 25616 3229 25636 3263
rect 25562 3153 25636 3229
rect 25692 3220 25703 3272
rect 25755 3220 25766 3272
rect 26082 3272 26156 3279
rect 25692 3213 25766 3220
rect 25822 3263 25896 3269
rect 25822 3229 25842 3263
rect 25876 3229 25896 3263
rect 25822 3153 25896 3229
rect 25952 3263 26026 3269
rect 25952 3229 25972 3263
rect 26006 3229 26026 3263
rect 25952 3153 26026 3229
rect 26082 3220 26093 3272
rect 26145 3220 26156 3272
rect 26472 3272 26546 3279
rect 26082 3213 26156 3220
rect 26212 3263 26286 3269
rect 26212 3229 26232 3263
rect 26266 3229 26286 3263
rect 26212 3153 26286 3229
rect 26342 3263 26416 3269
rect 26342 3229 26362 3263
rect 26396 3229 26416 3263
rect 26342 3153 26416 3229
rect 26472 3220 26483 3272
rect 26535 3220 26546 3272
rect 26472 3213 26546 3220
rect 26602 3263 26676 3269
rect 26602 3229 26622 3263
rect 26656 3229 26676 3263
rect 26602 3153 26676 3229
rect 12998 3139 15502 3153
rect 12998 3130 13267 3139
rect 12998 3096 13022 3130
rect 13056 3096 13104 3130
rect 13138 3096 13196 3130
rect 13230 3096 13267 3130
rect 12998 3087 13267 3096
rect 13319 3087 13331 3139
rect 13383 3087 13395 3139
rect 13447 3130 14047 3139
rect 13447 3096 13484 3130
rect 13518 3096 13586 3130
rect 13620 3096 13658 3130
rect 13692 3096 13730 3130
rect 13764 3096 13802 3130
rect 13836 3096 13874 3130
rect 13908 3096 13976 3130
rect 14010 3096 14047 3130
rect 13447 3087 14047 3096
rect 14099 3087 14111 3139
rect 14163 3087 14175 3139
rect 14227 3130 14827 3139
rect 14227 3096 14264 3130
rect 14298 3096 14366 3130
rect 14400 3096 14438 3130
rect 14472 3096 14510 3130
rect 14544 3096 14582 3130
rect 14616 3096 14654 3130
rect 14688 3096 14756 3130
rect 14790 3096 14827 3130
rect 14227 3087 14827 3096
rect 14879 3087 14891 3139
rect 14943 3087 14955 3139
rect 15007 3130 15502 3139
rect 15007 3096 15044 3130
rect 15078 3096 15146 3130
rect 15180 3096 15218 3130
rect 15252 3096 15290 3130
rect 15324 3096 15362 3130
rect 15396 3096 15434 3130
rect 15468 3096 15502 3130
rect 15007 3087 15502 3096
rect 12998 3073 15502 3087
rect 24590 3139 27094 3153
rect 24590 3130 24859 3139
rect 24590 3096 24614 3130
rect 24648 3096 24696 3130
rect 24730 3096 24788 3130
rect 24822 3096 24859 3130
rect 24590 3087 24859 3096
rect 24911 3087 24923 3139
rect 24975 3087 24987 3139
rect 25039 3130 25639 3139
rect 25039 3096 25076 3130
rect 25110 3096 25178 3130
rect 25212 3096 25250 3130
rect 25284 3096 25322 3130
rect 25356 3096 25394 3130
rect 25428 3096 25466 3130
rect 25500 3096 25568 3130
rect 25602 3096 25639 3130
rect 25039 3087 25639 3096
rect 25691 3087 25703 3139
rect 25755 3087 25767 3139
rect 25819 3130 26419 3139
rect 25819 3096 25856 3130
rect 25890 3096 25958 3130
rect 25992 3096 26030 3130
rect 26064 3096 26102 3130
rect 26136 3096 26174 3130
rect 26208 3096 26246 3130
rect 26280 3096 26348 3130
rect 26382 3096 26419 3130
rect 25819 3087 26419 3096
rect 26471 3087 26483 3139
rect 26535 3087 26547 3139
rect 26599 3130 27094 3139
rect 26599 3096 26636 3130
rect 26670 3096 26738 3130
rect 26772 3096 26810 3130
rect 26844 3096 26882 3130
rect 26916 3096 26954 3130
rect 26988 3096 27026 3130
rect 27060 3096 27094 3130
rect 26599 3087 27094 3096
rect 24590 3073 27094 3087
rect 12677 3006 12751 3013
rect 12677 2954 12688 3006
rect 12740 2954 12751 3006
rect 13190 2997 13264 3073
rect 13190 2963 13210 2997
rect 13244 2963 13264 2997
rect 13190 2957 13264 2963
rect 13320 3006 13394 3013
rect 12677 2947 12751 2954
rect 13320 2954 13331 3006
rect 13383 2954 13394 3006
rect 13450 2997 13524 3073
rect 13450 2963 13470 2997
rect 13504 2963 13524 2997
rect 13450 2957 13524 2963
rect 13580 2997 13654 3073
rect 13580 2963 13600 2997
rect 13634 2963 13654 2997
rect 13580 2957 13654 2963
rect 13710 3006 13784 3013
rect 13320 2947 13394 2954
rect 13710 2954 13721 3006
rect 13773 2954 13784 3006
rect 13840 2997 13914 3073
rect 13840 2963 13860 2997
rect 13894 2963 13914 2997
rect 13840 2957 13914 2963
rect 13970 2997 14044 3073
rect 13970 2963 13990 2997
rect 14024 2963 14044 2997
rect 13970 2957 14044 2963
rect 14100 3006 14174 3013
rect 13710 2947 13784 2954
rect 14100 2954 14111 3006
rect 14163 2954 14174 3006
rect 14230 2997 14304 3073
rect 14230 2963 14250 2997
rect 14284 2963 14304 2997
rect 14230 2957 14304 2963
rect 14360 2997 14434 3073
rect 14360 2963 14380 2997
rect 14414 2963 14434 2997
rect 14360 2957 14434 2963
rect 14490 3006 14564 3013
rect 14100 2947 14174 2954
rect 14490 2954 14501 3006
rect 14553 2954 14564 3006
rect 14620 2997 14694 3073
rect 14620 2963 14640 2997
rect 14674 2963 14694 2997
rect 14620 2957 14694 2963
rect 14750 2997 14824 3073
rect 14750 2963 14770 2997
rect 14804 2963 14824 2997
rect 14750 2957 14824 2963
rect 14880 3006 14954 3013
rect 14490 2947 14564 2954
rect 14880 2954 14891 3006
rect 14943 2954 14954 3006
rect 15010 2997 15084 3073
rect 15010 2963 15030 2997
rect 15064 2963 15084 2997
rect 15010 2957 15084 2963
rect 15140 2997 15214 3073
rect 15140 2963 15160 2997
rect 15194 2963 15214 2997
rect 15140 2957 15214 2963
rect 15270 3006 15344 3013
rect 14880 2947 14954 2954
rect 15270 2954 15281 3006
rect 15333 2954 15344 3006
rect 15400 2997 15474 3073
rect 15400 2963 15420 2997
rect 15454 2963 15474 2997
rect 15400 2957 15474 2963
rect 24269 3006 24343 3013
rect 15270 2947 15344 2954
rect 24269 2954 24280 3006
rect 24332 2954 24343 3006
rect 24782 2997 24856 3073
rect 24782 2963 24802 2997
rect 24836 2963 24856 2997
rect 24782 2957 24856 2963
rect 24912 3006 24986 3013
rect 24269 2947 24343 2954
rect 24912 2954 24923 3006
rect 24975 2954 24986 3006
rect 25042 2997 25116 3073
rect 25042 2963 25062 2997
rect 25096 2963 25116 2997
rect 25042 2957 25116 2963
rect 25172 2997 25246 3073
rect 25172 2963 25192 2997
rect 25226 2963 25246 2997
rect 25172 2957 25246 2963
rect 25302 3006 25376 3013
rect 24912 2947 24986 2954
rect 25302 2954 25313 3006
rect 25365 2954 25376 3006
rect 25432 2997 25506 3073
rect 25432 2963 25452 2997
rect 25486 2963 25506 2997
rect 25432 2957 25506 2963
rect 25562 2997 25636 3073
rect 25562 2963 25582 2997
rect 25616 2963 25636 2997
rect 25562 2957 25636 2963
rect 25692 3006 25766 3013
rect 25302 2947 25376 2954
rect 25692 2954 25703 3006
rect 25755 2954 25766 3006
rect 25822 2997 25896 3073
rect 25822 2963 25842 2997
rect 25876 2963 25896 2997
rect 25822 2957 25896 2963
rect 25952 2997 26026 3073
rect 25952 2963 25972 2997
rect 26006 2963 26026 2997
rect 25952 2957 26026 2963
rect 26082 3006 26156 3013
rect 25692 2947 25766 2954
rect 26082 2954 26093 3006
rect 26145 2954 26156 3006
rect 26212 2997 26286 3073
rect 26212 2963 26232 2997
rect 26266 2963 26286 2997
rect 26212 2957 26286 2963
rect 26342 2997 26416 3073
rect 26342 2963 26362 2997
rect 26396 2963 26416 2997
rect 26342 2957 26416 2963
rect 26472 3006 26546 3013
rect 26082 2947 26156 2954
rect 26472 2954 26483 3006
rect 26535 2954 26546 3006
rect 26602 2997 26676 3073
rect 26602 2963 26622 2997
rect 26656 2963 26676 2997
rect 26602 2957 26676 2963
rect 26732 2997 26806 3073
rect 26732 2963 26752 2997
rect 26786 2963 26806 2997
rect 26732 2957 26806 2963
rect 26862 3006 26936 3013
rect 26472 2947 26546 2954
rect 26862 2954 26873 3006
rect 26925 2954 26936 3006
rect 26992 2997 27066 3073
rect 26992 2963 27012 2997
rect 27046 2963 27066 2997
rect 26992 2957 27066 2963
rect 26862 2947 26936 2954
rect 13139 2860 13185 2872
rect 13139 2857 13145 2860
rect 13125 2833 13145 2857
rect 13179 2857 13185 2860
rect 13269 2860 13315 2872
rect 13269 2857 13275 2860
rect 13179 2833 13199 2857
rect 13125 2781 13136 2833
rect 13188 2781 13199 2833
rect 13125 2757 13145 2781
rect 13139 2754 13145 2757
rect 13179 2757 13199 2781
rect 13255 2833 13275 2857
rect 13309 2857 13315 2860
rect 13399 2860 13445 2872
rect 13309 2833 13329 2857
rect 13255 2781 13266 2833
rect 13318 2781 13329 2833
rect 13255 2757 13275 2781
rect 13179 2754 13185 2757
rect 13139 2742 13185 2754
rect 13269 2754 13275 2757
rect 13309 2757 13329 2781
rect 13399 2826 13405 2860
rect 13439 2826 13445 2860
rect 13529 2860 13575 2872
rect 13529 2857 13535 2860
rect 13399 2788 13445 2826
rect 13309 2754 13315 2757
rect 13269 2742 13315 2754
rect 13399 2754 13405 2788
rect 13439 2754 13445 2788
rect 13515 2833 13535 2857
rect 13569 2857 13575 2860
rect 13659 2860 13705 2872
rect 13659 2857 13665 2860
rect 13569 2833 13589 2857
rect 13515 2781 13526 2833
rect 13578 2781 13589 2833
rect 13515 2757 13535 2781
rect 13130 2517 13194 2524
rect 13130 2465 13136 2517
rect 13188 2465 13194 2517
rect 13130 2453 13194 2465
rect 13130 2401 13136 2453
rect 13188 2401 13194 2453
rect 13130 2394 13194 2401
rect 13260 2517 13324 2524
rect 13260 2465 13266 2517
rect 13318 2465 13324 2517
rect 13260 2453 13324 2465
rect 13260 2401 13266 2453
rect 13318 2401 13324 2453
rect 13260 2394 13324 2401
rect 13399 2512 13445 2754
rect 13529 2754 13535 2757
rect 13569 2757 13589 2781
rect 13645 2833 13665 2857
rect 13699 2857 13705 2860
rect 13789 2860 13835 2872
rect 13699 2833 13719 2857
rect 13645 2781 13656 2833
rect 13708 2781 13719 2833
rect 13645 2757 13665 2781
rect 13569 2754 13575 2757
rect 13529 2742 13575 2754
rect 13659 2754 13665 2757
rect 13699 2757 13719 2781
rect 13789 2826 13795 2860
rect 13829 2826 13835 2860
rect 13919 2860 13965 2872
rect 13919 2857 13925 2860
rect 13789 2788 13835 2826
rect 13699 2754 13705 2757
rect 13659 2742 13705 2754
rect 13789 2754 13795 2788
rect 13829 2754 13835 2788
rect 13905 2833 13925 2857
rect 13959 2857 13965 2860
rect 14049 2860 14095 2872
rect 14049 2857 14055 2860
rect 13959 2833 13979 2857
rect 13905 2781 13916 2833
rect 13968 2781 13979 2833
rect 13905 2757 13925 2781
rect 13399 2478 13405 2512
rect 13439 2478 13445 2512
rect 13399 2440 13445 2478
rect 13399 2406 13405 2440
rect 13439 2406 13445 2440
rect 13399 2394 13445 2406
rect 13520 2517 13584 2524
rect 13520 2465 13526 2517
rect 13578 2465 13584 2517
rect 13520 2453 13584 2465
rect 13520 2401 13526 2453
rect 13578 2401 13584 2453
rect 13520 2394 13584 2401
rect 13650 2517 13714 2524
rect 13650 2465 13656 2517
rect 13708 2465 13714 2517
rect 13650 2453 13714 2465
rect 13650 2401 13656 2453
rect 13708 2401 13714 2453
rect 13650 2394 13714 2401
rect 13789 2512 13835 2754
rect 13919 2754 13925 2757
rect 13959 2757 13979 2781
rect 14035 2833 14055 2857
rect 14089 2857 14095 2860
rect 14179 2860 14225 2872
rect 14089 2833 14109 2857
rect 14035 2781 14046 2833
rect 14098 2781 14109 2833
rect 14035 2757 14055 2781
rect 13959 2754 13965 2757
rect 13919 2742 13965 2754
rect 14049 2754 14055 2757
rect 14089 2757 14109 2781
rect 14179 2826 14185 2860
rect 14219 2826 14225 2860
rect 14309 2860 14355 2872
rect 14309 2857 14315 2860
rect 14179 2788 14225 2826
rect 14089 2754 14095 2757
rect 14049 2742 14095 2754
rect 14179 2754 14185 2788
rect 14219 2754 14225 2788
rect 14295 2833 14315 2857
rect 14349 2857 14355 2860
rect 14439 2860 14485 2872
rect 14439 2857 14445 2860
rect 14349 2833 14369 2857
rect 14295 2781 14306 2833
rect 14358 2781 14369 2833
rect 14295 2757 14315 2781
rect 13789 2478 13795 2512
rect 13829 2478 13835 2512
rect 13789 2440 13835 2478
rect 13789 2406 13795 2440
rect 13829 2406 13835 2440
rect 13789 2394 13835 2406
rect 13910 2517 13974 2524
rect 13910 2465 13916 2517
rect 13968 2465 13974 2517
rect 13910 2453 13974 2465
rect 13910 2401 13916 2453
rect 13968 2401 13974 2453
rect 13910 2394 13974 2401
rect 14040 2517 14104 2524
rect 14040 2465 14046 2517
rect 14098 2465 14104 2517
rect 14040 2453 14104 2465
rect 14040 2401 14046 2453
rect 14098 2401 14104 2453
rect 14040 2394 14104 2401
rect 14179 2512 14225 2754
rect 14309 2754 14315 2757
rect 14349 2757 14369 2781
rect 14425 2833 14445 2857
rect 14479 2857 14485 2860
rect 14569 2860 14615 2872
rect 14479 2833 14499 2857
rect 14425 2781 14436 2833
rect 14488 2781 14499 2833
rect 14425 2757 14445 2781
rect 14349 2754 14355 2757
rect 14309 2742 14355 2754
rect 14439 2754 14445 2757
rect 14479 2757 14499 2781
rect 14569 2826 14575 2860
rect 14609 2826 14615 2860
rect 14699 2860 14745 2872
rect 14699 2857 14705 2860
rect 14569 2788 14615 2826
rect 14479 2754 14485 2757
rect 14439 2742 14485 2754
rect 14569 2754 14575 2788
rect 14609 2754 14615 2788
rect 14685 2833 14705 2857
rect 14739 2857 14745 2860
rect 14829 2860 14875 2872
rect 14829 2857 14835 2860
rect 14739 2833 14759 2857
rect 14685 2781 14696 2833
rect 14748 2781 14759 2833
rect 14685 2757 14705 2781
rect 14179 2478 14185 2512
rect 14219 2478 14225 2512
rect 14179 2440 14225 2478
rect 14179 2406 14185 2440
rect 14219 2406 14225 2440
rect 14179 2394 14225 2406
rect 14300 2517 14364 2524
rect 14300 2465 14306 2517
rect 14358 2465 14364 2517
rect 14300 2453 14364 2465
rect 14300 2401 14306 2453
rect 14358 2401 14364 2453
rect 14300 2394 14364 2401
rect 14430 2517 14494 2524
rect 14430 2465 14436 2517
rect 14488 2465 14494 2517
rect 14430 2453 14494 2465
rect 14430 2401 14436 2453
rect 14488 2401 14494 2453
rect 14430 2394 14494 2401
rect 14569 2512 14615 2754
rect 14699 2754 14705 2757
rect 14739 2757 14759 2781
rect 14815 2833 14835 2857
rect 14869 2857 14875 2860
rect 14959 2860 15005 2872
rect 14869 2833 14889 2857
rect 14815 2781 14826 2833
rect 14878 2781 14889 2833
rect 14815 2757 14835 2781
rect 14739 2754 14745 2757
rect 14699 2742 14745 2754
rect 14829 2754 14835 2757
rect 14869 2757 14889 2781
rect 14959 2826 14965 2860
rect 14999 2826 15005 2860
rect 15089 2860 15135 2872
rect 15089 2857 15095 2860
rect 14959 2788 15005 2826
rect 14869 2754 14875 2757
rect 14829 2742 14875 2754
rect 14959 2754 14965 2788
rect 14999 2754 15005 2788
rect 15075 2833 15095 2857
rect 15129 2857 15135 2860
rect 15219 2860 15265 2872
rect 15219 2857 15225 2860
rect 15129 2833 15149 2857
rect 15075 2781 15086 2833
rect 15138 2781 15149 2833
rect 15075 2757 15095 2781
rect 14569 2478 14575 2512
rect 14609 2478 14615 2512
rect 14569 2440 14615 2478
rect 14569 2406 14575 2440
rect 14609 2406 14615 2440
rect 14569 2394 14615 2406
rect 14690 2517 14754 2524
rect 14690 2465 14696 2517
rect 14748 2465 14754 2517
rect 14690 2453 14754 2465
rect 14690 2401 14696 2453
rect 14748 2401 14754 2453
rect 14690 2394 14754 2401
rect 14820 2517 14884 2524
rect 14820 2465 14826 2517
rect 14878 2465 14884 2517
rect 14820 2453 14884 2465
rect 14820 2401 14826 2453
rect 14878 2401 14884 2453
rect 14820 2394 14884 2401
rect 14959 2512 15005 2754
rect 15089 2754 15095 2757
rect 15129 2757 15149 2781
rect 15205 2833 15225 2857
rect 15259 2857 15265 2860
rect 15349 2860 15395 2872
rect 15259 2833 15279 2857
rect 15205 2781 15216 2833
rect 15268 2781 15279 2833
rect 15205 2757 15225 2781
rect 15129 2754 15135 2757
rect 15089 2742 15135 2754
rect 15219 2754 15225 2757
rect 15259 2757 15279 2781
rect 15349 2826 15355 2860
rect 15389 2826 15395 2860
rect 15479 2860 15525 2872
rect 15479 2857 15485 2860
rect 15349 2788 15395 2826
rect 15259 2754 15265 2757
rect 15219 2742 15265 2754
rect 15349 2754 15355 2788
rect 15389 2754 15395 2788
rect 15465 2833 15485 2857
rect 15519 2857 15525 2860
rect 24731 2860 24777 2872
rect 24731 2857 24737 2860
rect 15519 2833 15539 2857
rect 15465 2781 15476 2833
rect 15528 2781 15539 2833
rect 15465 2757 15485 2781
rect 14959 2478 14965 2512
rect 14999 2478 15005 2512
rect 14959 2440 15005 2478
rect 14959 2406 14965 2440
rect 14999 2406 15005 2440
rect 14959 2394 15005 2406
rect 15080 2517 15144 2524
rect 15080 2465 15086 2517
rect 15138 2465 15144 2517
rect 15080 2453 15144 2465
rect 15080 2401 15086 2453
rect 15138 2401 15144 2453
rect 15080 2394 15144 2401
rect 15210 2517 15274 2524
rect 15210 2465 15216 2517
rect 15268 2465 15274 2517
rect 15210 2453 15274 2465
rect 15210 2401 15216 2453
rect 15268 2401 15274 2453
rect 15210 2394 15274 2401
rect 15349 2512 15395 2754
rect 15479 2754 15485 2757
rect 15519 2757 15539 2781
rect 24717 2833 24737 2857
rect 24771 2857 24777 2860
rect 24861 2860 24907 2872
rect 24861 2857 24867 2860
rect 24771 2833 24791 2857
rect 24717 2781 24728 2833
rect 24780 2781 24791 2833
rect 24717 2757 24737 2781
rect 15519 2754 15525 2757
rect 15479 2742 15525 2754
rect 24731 2754 24737 2757
rect 24771 2757 24791 2781
rect 24847 2833 24867 2857
rect 24901 2857 24907 2860
rect 24991 2860 25037 2872
rect 24901 2833 24921 2857
rect 24847 2781 24858 2833
rect 24910 2781 24921 2833
rect 24847 2757 24867 2781
rect 24771 2754 24777 2757
rect 24731 2742 24777 2754
rect 24861 2754 24867 2757
rect 24901 2757 24921 2781
rect 24991 2826 24997 2860
rect 25031 2826 25037 2860
rect 25121 2860 25167 2872
rect 25121 2857 25127 2860
rect 24991 2788 25037 2826
rect 24901 2754 24907 2757
rect 24861 2742 24907 2754
rect 24991 2754 24997 2788
rect 25031 2754 25037 2788
rect 25107 2833 25127 2857
rect 25161 2857 25167 2860
rect 25251 2860 25297 2872
rect 25251 2857 25257 2860
rect 25161 2833 25181 2857
rect 25107 2781 25118 2833
rect 25170 2781 25181 2833
rect 25107 2757 25127 2781
rect 15349 2478 15355 2512
rect 15389 2478 15395 2512
rect 15349 2440 15395 2478
rect 15349 2406 15355 2440
rect 15389 2406 15395 2440
rect 15349 2394 15395 2406
rect 24722 2517 24786 2524
rect 24722 2465 24728 2517
rect 24780 2465 24786 2517
rect 24722 2453 24786 2465
rect 24722 2401 24728 2453
rect 24780 2401 24786 2453
rect 24722 2394 24786 2401
rect 24852 2517 24916 2524
rect 24852 2465 24858 2517
rect 24910 2465 24916 2517
rect 24852 2453 24916 2465
rect 24852 2401 24858 2453
rect 24910 2401 24916 2453
rect 24852 2394 24916 2401
rect 24991 2512 25037 2754
rect 25121 2754 25127 2757
rect 25161 2757 25181 2781
rect 25237 2833 25257 2857
rect 25291 2857 25297 2860
rect 25381 2860 25427 2872
rect 25291 2833 25311 2857
rect 25237 2781 25248 2833
rect 25300 2781 25311 2833
rect 25237 2757 25257 2781
rect 25161 2754 25167 2757
rect 25121 2742 25167 2754
rect 25251 2754 25257 2757
rect 25291 2757 25311 2781
rect 25381 2826 25387 2860
rect 25421 2826 25427 2860
rect 25511 2860 25557 2872
rect 25511 2857 25517 2860
rect 25381 2788 25427 2826
rect 25291 2754 25297 2757
rect 25251 2742 25297 2754
rect 25381 2754 25387 2788
rect 25421 2754 25427 2788
rect 25497 2833 25517 2857
rect 25551 2857 25557 2860
rect 25641 2860 25687 2872
rect 25641 2857 25647 2860
rect 25551 2833 25571 2857
rect 25497 2781 25508 2833
rect 25560 2781 25571 2833
rect 25497 2757 25517 2781
rect 24991 2478 24997 2512
rect 25031 2478 25037 2512
rect 24991 2440 25037 2478
rect 24991 2406 24997 2440
rect 25031 2406 25037 2440
rect 24991 2394 25037 2406
rect 25112 2517 25176 2524
rect 25112 2465 25118 2517
rect 25170 2465 25176 2517
rect 25112 2453 25176 2465
rect 25112 2401 25118 2453
rect 25170 2401 25176 2453
rect 25112 2394 25176 2401
rect 25242 2517 25306 2524
rect 25242 2465 25248 2517
rect 25300 2465 25306 2517
rect 25242 2453 25306 2465
rect 25242 2401 25248 2453
rect 25300 2401 25306 2453
rect 25242 2394 25306 2401
rect 25381 2512 25427 2754
rect 25511 2754 25517 2757
rect 25551 2757 25571 2781
rect 25627 2833 25647 2857
rect 25681 2857 25687 2860
rect 25771 2860 25817 2872
rect 25681 2833 25701 2857
rect 25627 2781 25638 2833
rect 25690 2781 25701 2833
rect 25627 2757 25647 2781
rect 25551 2754 25557 2757
rect 25511 2742 25557 2754
rect 25641 2754 25647 2757
rect 25681 2757 25701 2781
rect 25771 2826 25777 2860
rect 25811 2826 25817 2860
rect 25901 2860 25947 2872
rect 25901 2857 25907 2860
rect 25771 2788 25817 2826
rect 25681 2754 25687 2757
rect 25641 2742 25687 2754
rect 25771 2754 25777 2788
rect 25811 2754 25817 2788
rect 25887 2833 25907 2857
rect 25941 2857 25947 2860
rect 26031 2860 26077 2872
rect 26031 2857 26037 2860
rect 25941 2833 25961 2857
rect 25887 2781 25898 2833
rect 25950 2781 25961 2833
rect 25887 2757 25907 2781
rect 25381 2478 25387 2512
rect 25421 2478 25427 2512
rect 25381 2440 25427 2478
rect 25381 2406 25387 2440
rect 25421 2406 25427 2440
rect 25381 2394 25427 2406
rect 25502 2517 25566 2524
rect 25502 2465 25508 2517
rect 25560 2465 25566 2517
rect 25502 2453 25566 2465
rect 25502 2401 25508 2453
rect 25560 2401 25566 2453
rect 25502 2394 25566 2401
rect 25632 2517 25696 2524
rect 25632 2465 25638 2517
rect 25690 2465 25696 2517
rect 25632 2453 25696 2465
rect 25632 2401 25638 2453
rect 25690 2401 25696 2453
rect 25632 2394 25696 2401
rect 25771 2512 25817 2754
rect 25901 2754 25907 2757
rect 25941 2757 25961 2781
rect 26017 2833 26037 2857
rect 26071 2857 26077 2860
rect 26161 2860 26207 2872
rect 26071 2833 26091 2857
rect 26017 2781 26028 2833
rect 26080 2781 26091 2833
rect 26017 2757 26037 2781
rect 25941 2754 25947 2757
rect 25901 2742 25947 2754
rect 26031 2754 26037 2757
rect 26071 2757 26091 2781
rect 26161 2826 26167 2860
rect 26201 2826 26207 2860
rect 26291 2860 26337 2872
rect 26291 2857 26297 2860
rect 26161 2788 26207 2826
rect 26071 2754 26077 2757
rect 26031 2742 26077 2754
rect 26161 2754 26167 2788
rect 26201 2754 26207 2788
rect 26277 2833 26297 2857
rect 26331 2857 26337 2860
rect 26421 2860 26467 2872
rect 26421 2857 26427 2860
rect 26331 2833 26351 2857
rect 26277 2781 26288 2833
rect 26340 2781 26351 2833
rect 26277 2757 26297 2781
rect 25771 2478 25777 2512
rect 25811 2478 25817 2512
rect 25771 2440 25817 2478
rect 25771 2406 25777 2440
rect 25811 2406 25817 2440
rect 25771 2394 25817 2406
rect 25892 2517 25956 2524
rect 25892 2465 25898 2517
rect 25950 2465 25956 2517
rect 25892 2453 25956 2465
rect 25892 2401 25898 2453
rect 25950 2401 25956 2453
rect 25892 2394 25956 2401
rect 26022 2517 26086 2524
rect 26022 2465 26028 2517
rect 26080 2465 26086 2517
rect 26022 2453 26086 2465
rect 26022 2401 26028 2453
rect 26080 2401 26086 2453
rect 26022 2394 26086 2401
rect 26161 2512 26207 2754
rect 26291 2754 26297 2757
rect 26331 2757 26351 2781
rect 26407 2833 26427 2857
rect 26461 2857 26467 2860
rect 26551 2860 26597 2872
rect 26461 2833 26481 2857
rect 26407 2781 26418 2833
rect 26470 2781 26481 2833
rect 26407 2757 26427 2781
rect 26331 2754 26337 2757
rect 26291 2742 26337 2754
rect 26421 2754 26427 2757
rect 26461 2757 26481 2781
rect 26551 2826 26557 2860
rect 26591 2826 26597 2860
rect 26681 2860 26727 2872
rect 26681 2857 26687 2860
rect 26551 2788 26597 2826
rect 26461 2754 26467 2757
rect 26421 2742 26467 2754
rect 26551 2754 26557 2788
rect 26591 2754 26597 2788
rect 26667 2833 26687 2857
rect 26721 2857 26727 2860
rect 26811 2860 26857 2872
rect 26811 2857 26817 2860
rect 26721 2833 26741 2857
rect 26667 2781 26678 2833
rect 26730 2781 26741 2833
rect 26667 2757 26687 2781
rect 26161 2478 26167 2512
rect 26201 2478 26207 2512
rect 26161 2440 26207 2478
rect 26161 2406 26167 2440
rect 26201 2406 26207 2440
rect 26161 2394 26207 2406
rect 26282 2517 26346 2524
rect 26282 2465 26288 2517
rect 26340 2465 26346 2517
rect 26282 2453 26346 2465
rect 26282 2401 26288 2453
rect 26340 2401 26346 2453
rect 26282 2394 26346 2401
rect 26412 2517 26476 2524
rect 26412 2465 26418 2517
rect 26470 2465 26476 2517
rect 26412 2453 26476 2465
rect 26412 2401 26418 2453
rect 26470 2401 26476 2453
rect 26412 2394 26476 2401
rect 26551 2512 26597 2754
rect 26681 2754 26687 2757
rect 26721 2757 26741 2781
rect 26797 2833 26817 2857
rect 26851 2857 26857 2860
rect 26941 2860 26987 2872
rect 26851 2833 26871 2857
rect 26797 2781 26808 2833
rect 26860 2781 26871 2833
rect 26797 2757 26817 2781
rect 26721 2754 26727 2757
rect 26681 2742 26727 2754
rect 26811 2754 26817 2757
rect 26851 2757 26871 2781
rect 26941 2826 26947 2860
rect 26981 2826 26987 2860
rect 27071 2860 27117 2872
rect 27071 2857 27077 2860
rect 26941 2788 26987 2826
rect 26851 2754 26857 2757
rect 26811 2742 26857 2754
rect 26941 2754 26947 2788
rect 26981 2754 26987 2788
rect 27057 2833 27077 2857
rect 27111 2857 27117 2860
rect 27111 2833 27131 2857
rect 27057 2781 27068 2833
rect 27120 2781 27131 2833
rect 27057 2757 27077 2781
rect 26551 2478 26557 2512
rect 26591 2478 26597 2512
rect 26551 2440 26597 2478
rect 26551 2406 26557 2440
rect 26591 2406 26597 2440
rect 26551 2394 26597 2406
rect 26672 2517 26736 2524
rect 26672 2465 26678 2517
rect 26730 2465 26736 2517
rect 26672 2453 26736 2465
rect 26672 2401 26678 2453
rect 26730 2401 26736 2453
rect 26672 2394 26736 2401
rect 26802 2517 26866 2524
rect 26802 2465 26808 2517
rect 26860 2465 26866 2517
rect 26802 2453 26866 2465
rect 26802 2401 26808 2453
rect 26860 2401 26866 2453
rect 26802 2394 26866 2401
rect 26941 2512 26987 2754
rect 27071 2754 27077 2757
rect 27111 2757 27131 2781
rect 27111 2754 27117 2757
rect 27071 2742 27117 2754
rect 26941 2478 26947 2512
rect 26981 2478 26987 2512
rect 26941 2440 26987 2478
rect 26941 2406 26947 2440
rect 26981 2406 26987 2440
rect 26941 2394 26987 2406
rect 12499 2318 15729 2319
rect 12499 2266 12596 2318
rect 12648 2309 15729 2318
rect 12648 2275 13210 2309
rect 13244 2275 13600 2309
rect 13634 2275 14380 2309
rect 14414 2275 15160 2309
rect 15194 2275 15729 2309
rect 12648 2266 15729 2275
rect 12499 2265 15729 2266
rect 24091 2318 27321 2319
rect 24091 2266 24188 2318
rect 24240 2309 27321 2318
rect 24240 2275 24802 2309
rect 24836 2275 25192 2309
rect 25226 2275 25972 2309
rect 26006 2275 26752 2309
rect 26786 2275 27321 2309
rect 24240 2266 27321 2275
rect 24091 2265 27321 2266
rect 12891 2161 13324 2167
rect 12891 2109 12897 2161
rect 12949 2109 13266 2161
rect 13318 2109 13324 2161
rect 12891 2103 13324 2109
rect 13420 2161 13714 2167
rect 13420 2152 13656 2161
rect 13420 2118 13436 2152
rect 13470 2118 13656 2152
rect 13420 2109 13656 2118
rect 13708 2109 13714 2161
rect 13420 2103 13714 2109
rect 13810 2161 14104 2167
rect 13810 2152 14046 2161
rect 13810 2118 13826 2152
rect 13860 2118 14046 2152
rect 13810 2109 14046 2118
rect 14098 2109 14104 2161
rect 13810 2103 14104 2109
rect 14200 2161 14494 2167
rect 14200 2152 14436 2161
rect 14200 2118 14216 2152
rect 14250 2118 14436 2152
rect 14200 2109 14436 2118
rect 14488 2109 14494 2161
rect 14200 2103 14494 2109
rect 14590 2161 14884 2167
rect 14590 2152 14826 2161
rect 14590 2118 14606 2152
rect 14640 2118 14826 2152
rect 14590 2109 14826 2118
rect 14878 2109 14884 2161
rect 14590 2103 14884 2109
rect 14980 2161 15274 2167
rect 14980 2152 15216 2161
rect 14980 2118 14996 2152
rect 15030 2118 15216 2152
rect 14980 2109 15216 2118
rect 15268 2109 15274 2161
rect 14980 2103 15274 2109
rect 15370 2161 15729 2167
rect 15370 2152 15671 2161
rect 15370 2118 15386 2152
rect 15420 2118 15671 2152
rect 15370 2109 15671 2118
rect 15723 2109 15729 2161
rect 15370 2103 15729 2109
rect 24483 2161 24916 2167
rect 24483 2109 24489 2161
rect 24541 2109 24858 2161
rect 24910 2109 24916 2161
rect 24483 2103 24916 2109
rect 25012 2161 25306 2167
rect 25012 2152 25248 2161
rect 25012 2118 25028 2152
rect 25062 2118 25248 2152
rect 25012 2109 25248 2118
rect 25300 2109 25306 2161
rect 25012 2103 25306 2109
rect 25402 2161 25696 2167
rect 25402 2152 25638 2161
rect 25402 2118 25418 2152
rect 25452 2118 25638 2152
rect 25402 2109 25638 2118
rect 25690 2109 25696 2161
rect 25402 2103 25696 2109
rect 25792 2161 26086 2167
rect 25792 2152 26028 2161
rect 25792 2118 25808 2152
rect 25842 2118 26028 2152
rect 25792 2109 26028 2118
rect 26080 2109 26086 2161
rect 25792 2103 26086 2109
rect 26182 2161 26476 2167
rect 26182 2152 26418 2161
rect 26182 2118 26198 2152
rect 26232 2118 26418 2152
rect 26182 2109 26418 2118
rect 26470 2109 26476 2161
rect 26182 2103 26476 2109
rect 26572 2161 26866 2167
rect 26572 2152 26808 2161
rect 26572 2118 26588 2152
rect 26622 2118 26808 2152
rect 26572 2109 26808 2118
rect 26860 2109 26866 2161
rect 26572 2103 26866 2109
rect 26962 2161 27321 2167
rect 26962 2152 27263 2161
rect 26962 2118 26978 2152
rect 27012 2118 27263 2152
rect 26962 2109 27263 2118
rect 27315 2109 27321 2161
rect 26962 2103 27321 2109
rect 13260 1872 13324 1884
rect 13260 1865 13275 1872
rect 13309 1865 13324 1872
rect 13260 1813 13266 1865
rect 13318 1813 13324 1865
rect 13260 1801 13324 1813
rect 13260 1749 13266 1801
rect 13318 1749 13324 1801
rect 13260 1737 13324 1749
rect 13260 1685 13266 1737
rect 13318 1685 13324 1737
rect 13260 1673 13324 1685
rect 13260 1621 13266 1673
rect 13318 1621 13324 1673
rect 13260 1609 13324 1621
rect 13260 1557 13266 1609
rect 13318 1557 13324 1609
rect 13260 1550 13275 1557
rect 13309 1550 13324 1557
rect 13260 1538 13324 1550
rect 13399 1872 13445 1884
rect 13399 1838 13405 1872
rect 13439 1838 13445 1872
rect 13399 1800 13445 1838
rect 13399 1766 13405 1800
rect 13439 1766 13445 1800
rect 13399 1728 13445 1766
rect 13399 1694 13405 1728
rect 13439 1694 13445 1728
rect 13399 1656 13445 1694
rect 13399 1622 13405 1656
rect 13439 1622 13445 1656
rect 13399 1584 13445 1622
rect 13399 1550 13405 1584
rect 13439 1550 13445 1584
rect 13139 1324 13185 1336
rect 13139 1290 13145 1324
rect 13179 1290 13185 1324
rect 13139 1252 13185 1290
rect 13139 1218 13145 1252
rect 13179 1218 13185 1252
rect 13139 1213 13185 1218
rect 13269 1324 13315 1336
rect 13269 1290 13275 1324
rect 13309 1290 13315 1324
rect 13269 1252 13315 1290
rect 13269 1218 13275 1252
rect 13309 1218 13315 1252
rect 13269 1213 13315 1218
rect 13399 1324 13445 1550
rect 13650 1872 13714 1884
rect 13650 1865 13665 1872
rect 13699 1865 13714 1872
rect 13650 1813 13656 1865
rect 13708 1813 13714 1865
rect 13650 1801 13714 1813
rect 13650 1749 13656 1801
rect 13708 1749 13714 1801
rect 13650 1737 13714 1749
rect 13650 1685 13656 1737
rect 13708 1685 13714 1737
rect 13650 1673 13714 1685
rect 13650 1621 13656 1673
rect 13708 1621 13714 1673
rect 13650 1609 13714 1621
rect 13650 1557 13656 1609
rect 13708 1557 13714 1609
rect 13650 1550 13665 1557
rect 13699 1550 13714 1557
rect 13650 1538 13714 1550
rect 13789 1872 13835 1884
rect 13789 1838 13795 1872
rect 13829 1838 13835 1872
rect 13789 1800 13835 1838
rect 13789 1766 13795 1800
rect 13829 1766 13835 1800
rect 13789 1728 13835 1766
rect 13789 1694 13795 1728
rect 13829 1694 13835 1728
rect 13789 1656 13835 1694
rect 13789 1622 13795 1656
rect 13829 1622 13835 1656
rect 13789 1584 13835 1622
rect 13789 1550 13795 1584
rect 13829 1550 13835 1584
rect 13399 1290 13405 1324
rect 13439 1290 13445 1324
rect 13399 1252 13445 1290
rect 13399 1218 13405 1252
rect 13439 1218 13445 1252
rect 13125 1189 13199 1213
rect 13125 1137 13136 1189
rect 13188 1137 13199 1189
rect 13125 1113 13199 1137
rect 13255 1189 13329 1213
rect 13255 1137 13266 1189
rect 13318 1137 13329 1189
rect 13255 1113 13329 1137
rect 13399 1180 13445 1218
rect 13529 1324 13575 1336
rect 13529 1290 13535 1324
rect 13569 1290 13575 1324
rect 13529 1252 13575 1290
rect 13529 1218 13535 1252
rect 13569 1218 13575 1252
rect 13529 1213 13575 1218
rect 13659 1324 13705 1336
rect 13659 1290 13665 1324
rect 13699 1290 13705 1324
rect 13659 1252 13705 1290
rect 13659 1218 13665 1252
rect 13699 1218 13705 1252
rect 13659 1213 13705 1218
rect 13789 1324 13835 1550
rect 14040 1872 14104 1884
rect 14040 1865 14055 1872
rect 14089 1865 14104 1872
rect 14040 1813 14046 1865
rect 14098 1813 14104 1865
rect 14040 1801 14104 1813
rect 14040 1749 14046 1801
rect 14098 1749 14104 1801
rect 14040 1737 14104 1749
rect 14040 1685 14046 1737
rect 14098 1685 14104 1737
rect 14040 1673 14104 1685
rect 14040 1621 14046 1673
rect 14098 1621 14104 1673
rect 14040 1609 14104 1621
rect 14040 1557 14046 1609
rect 14098 1557 14104 1609
rect 14040 1550 14055 1557
rect 14089 1550 14104 1557
rect 14040 1538 14104 1550
rect 14179 1872 14225 1884
rect 14179 1838 14185 1872
rect 14219 1838 14225 1872
rect 14179 1800 14225 1838
rect 14179 1766 14185 1800
rect 14219 1766 14225 1800
rect 14179 1728 14225 1766
rect 14179 1694 14185 1728
rect 14219 1694 14225 1728
rect 14179 1656 14225 1694
rect 14179 1622 14185 1656
rect 14219 1622 14225 1656
rect 14179 1584 14225 1622
rect 14179 1550 14185 1584
rect 14219 1550 14225 1584
rect 13789 1290 13795 1324
rect 13829 1290 13835 1324
rect 13789 1252 13835 1290
rect 13789 1218 13795 1252
rect 13829 1218 13835 1252
rect 13399 1146 13405 1180
rect 13439 1146 13445 1180
rect 13139 1108 13185 1113
rect 13139 1074 13145 1108
rect 13179 1074 13185 1108
rect 13139 1036 13185 1074
rect 13139 1002 13145 1036
rect 13179 1002 13185 1036
rect 13139 990 13185 1002
rect 13269 1108 13315 1113
rect 13269 1074 13275 1108
rect 13309 1074 13315 1108
rect 13269 1036 13315 1074
rect 13269 1002 13275 1036
rect 13309 1002 13315 1036
rect 13269 990 13315 1002
rect 13399 1108 13445 1146
rect 13515 1189 13589 1213
rect 13515 1137 13526 1189
rect 13578 1137 13589 1189
rect 13515 1113 13589 1137
rect 13645 1189 13719 1213
rect 13645 1137 13656 1189
rect 13708 1137 13719 1189
rect 13645 1113 13719 1137
rect 13789 1180 13835 1218
rect 13919 1324 13965 1336
rect 13919 1290 13925 1324
rect 13959 1290 13965 1324
rect 13919 1252 13965 1290
rect 13919 1218 13925 1252
rect 13959 1218 13965 1252
rect 13919 1213 13965 1218
rect 14049 1324 14095 1336
rect 14049 1290 14055 1324
rect 14089 1290 14095 1324
rect 14049 1252 14095 1290
rect 14049 1218 14055 1252
rect 14089 1218 14095 1252
rect 14049 1213 14095 1218
rect 14179 1324 14225 1550
rect 14430 1872 14494 1884
rect 14430 1865 14445 1872
rect 14479 1865 14494 1872
rect 14430 1813 14436 1865
rect 14488 1813 14494 1865
rect 14430 1801 14494 1813
rect 14430 1749 14436 1801
rect 14488 1749 14494 1801
rect 14430 1737 14494 1749
rect 14430 1685 14436 1737
rect 14488 1685 14494 1737
rect 14430 1673 14494 1685
rect 14430 1621 14436 1673
rect 14488 1621 14494 1673
rect 14430 1609 14494 1621
rect 14430 1557 14436 1609
rect 14488 1557 14494 1609
rect 14430 1550 14445 1557
rect 14479 1550 14494 1557
rect 14430 1538 14494 1550
rect 14569 1872 14615 1884
rect 14569 1838 14575 1872
rect 14609 1838 14615 1872
rect 14569 1800 14615 1838
rect 14569 1766 14575 1800
rect 14609 1766 14615 1800
rect 14569 1728 14615 1766
rect 14569 1694 14575 1728
rect 14609 1694 14615 1728
rect 14569 1656 14615 1694
rect 14569 1622 14575 1656
rect 14609 1622 14615 1656
rect 14569 1584 14615 1622
rect 14569 1550 14575 1584
rect 14609 1550 14615 1584
rect 14179 1290 14185 1324
rect 14219 1290 14225 1324
rect 14179 1252 14225 1290
rect 14179 1218 14185 1252
rect 14219 1218 14225 1252
rect 13789 1146 13795 1180
rect 13829 1146 13835 1180
rect 13399 1074 13405 1108
rect 13439 1074 13445 1108
rect 13399 1036 13445 1074
rect 13399 1002 13405 1036
rect 13439 1002 13445 1036
rect 13399 990 13445 1002
rect 13529 1108 13575 1113
rect 13529 1074 13535 1108
rect 13569 1074 13575 1108
rect 13529 1036 13575 1074
rect 13529 1002 13535 1036
rect 13569 1002 13575 1036
rect 13529 990 13575 1002
rect 13659 1108 13705 1113
rect 13659 1074 13665 1108
rect 13699 1074 13705 1108
rect 13659 1036 13705 1074
rect 13659 1002 13665 1036
rect 13699 1002 13705 1036
rect 13659 990 13705 1002
rect 13789 1108 13835 1146
rect 13905 1189 13979 1213
rect 13905 1137 13916 1189
rect 13968 1137 13979 1189
rect 13905 1113 13979 1137
rect 14035 1189 14109 1213
rect 14035 1137 14046 1189
rect 14098 1137 14109 1189
rect 14035 1113 14109 1137
rect 14179 1180 14225 1218
rect 14309 1324 14355 1336
rect 14309 1290 14315 1324
rect 14349 1290 14355 1324
rect 14309 1252 14355 1290
rect 14309 1218 14315 1252
rect 14349 1218 14355 1252
rect 14309 1213 14355 1218
rect 14439 1324 14485 1336
rect 14439 1290 14445 1324
rect 14479 1290 14485 1324
rect 14439 1252 14485 1290
rect 14439 1218 14445 1252
rect 14479 1218 14485 1252
rect 14439 1213 14485 1218
rect 14569 1324 14615 1550
rect 14820 1872 14884 1884
rect 14820 1865 14835 1872
rect 14869 1865 14884 1872
rect 14820 1813 14826 1865
rect 14878 1813 14884 1865
rect 14820 1801 14884 1813
rect 14820 1749 14826 1801
rect 14878 1749 14884 1801
rect 14820 1737 14884 1749
rect 14820 1685 14826 1737
rect 14878 1685 14884 1737
rect 14820 1673 14884 1685
rect 14820 1621 14826 1673
rect 14878 1621 14884 1673
rect 14820 1609 14884 1621
rect 14820 1557 14826 1609
rect 14878 1557 14884 1609
rect 14820 1550 14835 1557
rect 14869 1550 14884 1557
rect 14820 1538 14884 1550
rect 14959 1872 15005 1884
rect 14959 1838 14965 1872
rect 14999 1838 15005 1872
rect 14959 1800 15005 1838
rect 14959 1766 14965 1800
rect 14999 1766 15005 1800
rect 14959 1728 15005 1766
rect 14959 1694 14965 1728
rect 14999 1694 15005 1728
rect 14959 1656 15005 1694
rect 14959 1622 14965 1656
rect 14999 1622 15005 1656
rect 14959 1584 15005 1622
rect 14959 1550 14965 1584
rect 14999 1550 15005 1584
rect 14569 1290 14575 1324
rect 14609 1290 14615 1324
rect 14569 1252 14615 1290
rect 14569 1218 14575 1252
rect 14609 1218 14615 1252
rect 14179 1146 14185 1180
rect 14219 1146 14225 1180
rect 13789 1074 13795 1108
rect 13829 1074 13835 1108
rect 13789 1036 13835 1074
rect 13789 1002 13795 1036
rect 13829 1002 13835 1036
rect 13789 990 13835 1002
rect 13919 1108 13965 1113
rect 13919 1074 13925 1108
rect 13959 1074 13965 1108
rect 13919 1036 13965 1074
rect 13919 1002 13925 1036
rect 13959 1002 13965 1036
rect 13919 990 13965 1002
rect 14049 1108 14095 1113
rect 14049 1074 14055 1108
rect 14089 1074 14095 1108
rect 14049 1036 14095 1074
rect 14049 1002 14055 1036
rect 14089 1002 14095 1036
rect 14049 990 14095 1002
rect 14179 1108 14225 1146
rect 14295 1189 14369 1213
rect 14295 1137 14306 1189
rect 14358 1137 14369 1189
rect 14295 1113 14369 1137
rect 14425 1189 14499 1213
rect 14425 1137 14436 1189
rect 14488 1137 14499 1189
rect 14425 1113 14499 1137
rect 14569 1180 14615 1218
rect 14699 1324 14745 1336
rect 14699 1290 14705 1324
rect 14739 1290 14745 1324
rect 14699 1252 14745 1290
rect 14699 1218 14705 1252
rect 14739 1218 14745 1252
rect 14699 1213 14745 1218
rect 14829 1324 14875 1336
rect 14829 1290 14835 1324
rect 14869 1290 14875 1324
rect 14829 1252 14875 1290
rect 14829 1218 14835 1252
rect 14869 1218 14875 1252
rect 14829 1213 14875 1218
rect 14959 1324 15005 1550
rect 15210 1872 15274 1884
rect 15210 1865 15225 1872
rect 15259 1865 15274 1872
rect 15210 1813 15216 1865
rect 15268 1813 15274 1865
rect 15210 1801 15274 1813
rect 15210 1749 15216 1801
rect 15268 1749 15274 1801
rect 15210 1737 15274 1749
rect 15210 1685 15216 1737
rect 15268 1685 15274 1737
rect 15210 1673 15274 1685
rect 15210 1621 15216 1673
rect 15268 1621 15274 1673
rect 15210 1609 15274 1621
rect 15210 1557 15216 1609
rect 15268 1557 15274 1609
rect 15210 1550 15225 1557
rect 15259 1550 15274 1557
rect 15210 1538 15274 1550
rect 15349 1872 15395 1884
rect 15349 1838 15355 1872
rect 15389 1838 15395 1872
rect 15349 1800 15395 1838
rect 15349 1766 15355 1800
rect 15389 1766 15395 1800
rect 15349 1728 15395 1766
rect 15349 1694 15355 1728
rect 15389 1694 15395 1728
rect 15349 1656 15395 1694
rect 15349 1622 15355 1656
rect 15389 1622 15395 1656
rect 15349 1584 15395 1622
rect 15349 1550 15355 1584
rect 15389 1550 15395 1584
rect 14959 1290 14965 1324
rect 14999 1290 15005 1324
rect 14959 1252 15005 1290
rect 14959 1218 14965 1252
rect 14999 1218 15005 1252
rect 14569 1146 14575 1180
rect 14609 1146 14615 1180
rect 14179 1074 14185 1108
rect 14219 1074 14225 1108
rect 14179 1036 14225 1074
rect 14179 1002 14185 1036
rect 14219 1002 14225 1036
rect 14179 990 14225 1002
rect 14309 1108 14355 1113
rect 14309 1074 14315 1108
rect 14349 1074 14355 1108
rect 14309 1036 14355 1074
rect 14309 1002 14315 1036
rect 14349 1002 14355 1036
rect 14309 990 14355 1002
rect 14439 1108 14485 1113
rect 14439 1074 14445 1108
rect 14479 1074 14485 1108
rect 14439 1036 14485 1074
rect 14439 1002 14445 1036
rect 14479 1002 14485 1036
rect 14439 990 14485 1002
rect 14569 1108 14615 1146
rect 14685 1189 14759 1213
rect 14685 1137 14696 1189
rect 14748 1137 14759 1189
rect 14685 1113 14759 1137
rect 14815 1189 14889 1213
rect 14815 1137 14826 1189
rect 14878 1137 14889 1189
rect 14815 1113 14889 1137
rect 14959 1180 15005 1218
rect 15089 1324 15135 1336
rect 15089 1290 15095 1324
rect 15129 1290 15135 1324
rect 15089 1252 15135 1290
rect 15089 1218 15095 1252
rect 15129 1218 15135 1252
rect 15089 1213 15135 1218
rect 15219 1324 15265 1336
rect 15219 1290 15225 1324
rect 15259 1290 15265 1324
rect 15219 1252 15265 1290
rect 15219 1218 15225 1252
rect 15259 1218 15265 1252
rect 15219 1213 15265 1218
rect 15349 1324 15395 1550
rect 24852 1872 24916 1884
rect 24852 1865 24867 1872
rect 24901 1865 24916 1872
rect 24852 1813 24858 1865
rect 24910 1813 24916 1865
rect 24852 1801 24916 1813
rect 24852 1749 24858 1801
rect 24910 1749 24916 1801
rect 24852 1737 24916 1749
rect 24852 1685 24858 1737
rect 24910 1685 24916 1737
rect 24852 1673 24916 1685
rect 24852 1621 24858 1673
rect 24910 1621 24916 1673
rect 24852 1609 24916 1621
rect 24852 1557 24858 1609
rect 24910 1557 24916 1609
rect 24852 1550 24867 1557
rect 24901 1550 24916 1557
rect 24852 1538 24916 1550
rect 24991 1872 25037 1884
rect 24991 1838 24997 1872
rect 25031 1838 25037 1872
rect 24991 1800 25037 1838
rect 24991 1766 24997 1800
rect 25031 1766 25037 1800
rect 24991 1728 25037 1766
rect 24991 1694 24997 1728
rect 25031 1694 25037 1728
rect 24991 1656 25037 1694
rect 24991 1622 24997 1656
rect 25031 1622 25037 1656
rect 24991 1584 25037 1622
rect 24991 1550 24997 1584
rect 25031 1550 25037 1584
rect 15349 1290 15355 1324
rect 15389 1290 15395 1324
rect 15349 1252 15395 1290
rect 15349 1218 15355 1252
rect 15389 1218 15395 1252
rect 14959 1146 14965 1180
rect 14999 1146 15005 1180
rect 14569 1074 14575 1108
rect 14609 1074 14615 1108
rect 14569 1036 14615 1074
rect 14569 1002 14575 1036
rect 14609 1002 14615 1036
rect 14569 990 14615 1002
rect 14699 1108 14745 1113
rect 14699 1074 14705 1108
rect 14739 1074 14745 1108
rect 14699 1036 14745 1074
rect 14699 1002 14705 1036
rect 14739 1002 14745 1036
rect 14699 990 14745 1002
rect 14829 1108 14875 1113
rect 14829 1074 14835 1108
rect 14869 1074 14875 1108
rect 14829 1036 14875 1074
rect 14829 1002 14835 1036
rect 14869 1002 14875 1036
rect 14829 990 14875 1002
rect 14959 1108 15005 1146
rect 15075 1189 15149 1213
rect 15075 1137 15086 1189
rect 15138 1137 15149 1189
rect 15075 1113 15149 1137
rect 15205 1189 15279 1213
rect 15205 1137 15216 1189
rect 15268 1137 15279 1189
rect 15205 1113 15279 1137
rect 15349 1180 15395 1218
rect 15479 1324 15525 1336
rect 15479 1290 15485 1324
rect 15519 1290 15525 1324
rect 15479 1252 15525 1290
rect 15479 1218 15485 1252
rect 15519 1218 15525 1252
rect 15479 1213 15525 1218
rect 24731 1324 24777 1336
rect 24731 1290 24737 1324
rect 24771 1290 24777 1324
rect 24731 1252 24777 1290
rect 24731 1218 24737 1252
rect 24771 1218 24777 1252
rect 24731 1213 24777 1218
rect 24861 1324 24907 1336
rect 24861 1290 24867 1324
rect 24901 1290 24907 1324
rect 24861 1252 24907 1290
rect 24861 1218 24867 1252
rect 24901 1218 24907 1252
rect 24861 1213 24907 1218
rect 24991 1324 25037 1550
rect 25242 1872 25306 1884
rect 25242 1865 25257 1872
rect 25291 1865 25306 1872
rect 25242 1813 25248 1865
rect 25300 1813 25306 1865
rect 25242 1801 25306 1813
rect 25242 1749 25248 1801
rect 25300 1749 25306 1801
rect 25242 1737 25306 1749
rect 25242 1685 25248 1737
rect 25300 1685 25306 1737
rect 25242 1673 25306 1685
rect 25242 1621 25248 1673
rect 25300 1621 25306 1673
rect 25242 1609 25306 1621
rect 25242 1557 25248 1609
rect 25300 1557 25306 1609
rect 25242 1550 25257 1557
rect 25291 1550 25306 1557
rect 25242 1538 25306 1550
rect 25381 1872 25427 1884
rect 25381 1838 25387 1872
rect 25421 1838 25427 1872
rect 25381 1800 25427 1838
rect 25381 1766 25387 1800
rect 25421 1766 25427 1800
rect 25381 1728 25427 1766
rect 25381 1694 25387 1728
rect 25421 1694 25427 1728
rect 25381 1656 25427 1694
rect 25381 1622 25387 1656
rect 25421 1622 25427 1656
rect 25381 1584 25427 1622
rect 25381 1550 25387 1584
rect 25421 1550 25427 1584
rect 24991 1290 24997 1324
rect 25031 1290 25037 1324
rect 24991 1252 25037 1290
rect 24991 1218 24997 1252
rect 25031 1218 25037 1252
rect 15349 1146 15355 1180
rect 15389 1146 15395 1180
rect 14959 1074 14965 1108
rect 14999 1074 15005 1108
rect 14959 1036 15005 1074
rect 14959 1002 14965 1036
rect 14999 1002 15005 1036
rect 14959 990 15005 1002
rect 15089 1108 15135 1113
rect 15089 1074 15095 1108
rect 15129 1074 15135 1108
rect 15089 1036 15135 1074
rect 15089 1002 15095 1036
rect 15129 1002 15135 1036
rect 15089 990 15135 1002
rect 15219 1108 15265 1113
rect 15219 1074 15225 1108
rect 15259 1074 15265 1108
rect 15219 1036 15265 1074
rect 15219 1002 15225 1036
rect 15259 1002 15265 1036
rect 15219 990 15265 1002
rect 15349 1108 15395 1146
rect 15465 1189 15539 1213
rect 15465 1137 15476 1189
rect 15528 1137 15539 1189
rect 15465 1113 15539 1137
rect 24717 1189 24791 1213
rect 24717 1137 24728 1189
rect 24780 1137 24791 1189
rect 24717 1113 24791 1137
rect 24847 1189 24921 1213
rect 24847 1137 24858 1189
rect 24910 1137 24921 1189
rect 24847 1113 24921 1137
rect 24991 1180 25037 1218
rect 25121 1324 25167 1336
rect 25121 1290 25127 1324
rect 25161 1290 25167 1324
rect 25121 1252 25167 1290
rect 25121 1218 25127 1252
rect 25161 1218 25167 1252
rect 25121 1213 25167 1218
rect 25251 1324 25297 1336
rect 25251 1290 25257 1324
rect 25291 1290 25297 1324
rect 25251 1252 25297 1290
rect 25251 1218 25257 1252
rect 25291 1218 25297 1252
rect 25251 1213 25297 1218
rect 25381 1324 25427 1550
rect 25632 1872 25696 1884
rect 25632 1865 25647 1872
rect 25681 1865 25696 1872
rect 25632 1813 25638 1865
rect 25690 1813 25696 1865
rect 25632 1801 25696 1813
rect 25632 1749 25638 1801
rect 25690 1749 25696 1801
rect 25632 1737 25696 1749
rect 25632 1685 25638 1737
rect 25690 1685 25696 1737
rect 25632 1673 25696 1685
rect 25632 1621 25638 1673
rect 25690 1621 25696 1673
rect 25632 1609 25696 1621
rect 25632 1557 25638 1609
rect 25690 1557 25696 1609
rect 25632 1550 25647 1557
rect 25681 1550 25696 1557
rect 25632 1538 25696 1550
rect 25771 1872 25817 1884
rect 25771 1838 25777 1872
rect 25811 1838 25817 1872
rect 25771 1800 25817 1838
rect 25771 1766 25777 1800
rect 25811 1766 25817 1800
rect 25771 1728 25817 1766
rect 25771 1694 25777 1728
rect 25811 1694 25817 1728
rect 25771 1656 25817 1694
rect 25771 1622 25777 1656
rect 25811 1622 25817 1656
rect 25771 1584 25817 1622
rect 25771 1550 25777 1584
rect 25811 1550 25817 1584
rect 25381 1290 25387 1324
rect 25421 1290 25427 1324
rect 25381 1252 25427 1290
rect 25381 1218 25387 1252
rect 25421 1218 25427 1252
rect 24991 1146 24997 1180
rect 25031 1146 25037 1180
rect 15349 1074 15355 1108
rect 15389 1074 15395 1108
rect 15349 1036 15395 1074
rect 15349 1002 15355 1036
rect 15389 1002 15395 1036
rect 15349 990 15395 1002
rect 15479 1108 15525 1113
rect 15479 1074 15485 1108
rect 15519 1074 15525 1108
rect 15479 1036 15525 1074
rect 15479 1002 15485 1036
rect 15519 1002 15525 1036
rect 15479 990 15525 1002
rect 24731 1108 24777 1113
rect 24731 1074 24737 1108
rect 24771 1074 24777 1108
rect 24731 1036 24777 1074
rect 24731 1002 24737 1036
rect 24771 1002 24777 1036
rect 24731 990 24777 1002
rect 24861 1108 24907 1113
rect 24861 1074 24867 1108
rect 24901 1074 24907 1108
rect 24861 1036 24907 1074
rect 24861 1002 24867 1036
rect 24901 1002 24907 1036
rect 24861 990 24907 1002
rect 24991 1108 25037 1146
rect 25107 1189 25181 1213
rect 25107 1137 25118 1189
rect 25170 1137 25181 1189
rect 25107 1113 25181 1137
rect 25237 1189 25311 1213
rect 25237 1137 25248 1189
rect 25300 1137 25311 1189
rect 25237 1113 25311 1137
rect 25381 1180 25427 1218
rect 25511 1324 25557 1336
rect 25511 1290 25517 1324
rect 25551 1290 25557 1324
rect 25511 1252 25557 1290
rect 25511 1218 25517 1252
rect 25551 1218 25557 1252
rect 25511 1213 25557 1218
rect 25641 1324 25687 1336
rect 25641 1290 25647 1324
rect 25681 1290 25687 1324
rect 25641 1252 25687 1290
rect 25641 1218 25647 1252
rect 25681 1218 25687 1252
rect 25641 1213 25687 1218
rect 25771 1324 25817 1550
rect 26022 1872 26086 1884
rect 26022 1865 26037 1872
rect 26071 1865 26086 1872
rect 26022 1813 26028 1865
rect 26080 1813 26086 1865
rect 26022 1801 26086 1813
rect 26022 1749 26028 1801
rect 26080 1749 26086 1801
rect 26022 1737 26086 1749
rect 26022 1685 26028 1737
rect 26080 1685 26086 1737
rect 26022 1673 26086 1685
rect 26022 1621 26028 1673
rect 26080 1621 26086 1673
rect 26022 1609 26086 1621
rect 26022 1557 26028 1609
rect 26080 1557 26086 1609
rect 26022 1550 26037 1557
rect 26071 1550 26086 1557
rect 26022 1538 26086 1550
rect 26161 1872 26207 1884
rect 26161 1838 26167 1872
rect 26201 1838 26207 1872
rect 26161 1800 26207 1838
rect 26161 1766 26167 1800
rect 26201 1766 26207 1800
rect 26161 1728 26207 1766
rect 26161 1694 26167 1728
rect 26201 1694 26207 1728
rect 26161 1656 26207 1694
rect 26161 1622 26167 1656
rect 26201 1622 26207 1656
rect 26161 1584 26207 1622
rect 26161 1550 26167 1584
rect 26201 1550 26207 1584
rect 25771 1290 25777 1324
rect 25811 1290 25817 1324
rect 25771 1252 25817 1290
rect 25771 1218 25777 1252
rect 25811 1218 25817 1252
rect 25381 1146 25387 1180
rect 25421 1146 25427 1180
rect 24991 1074 24997 1108
rect 25031 1074 25037 1108
rect 24991 1036 25037 1074
rect 24991 1002 24997 1036
rect 25031 1002 25037 1036
rect 24991 990 25037 1002
rect 25121 1108 25167 1113
rect 25121 1074 25127 1108
rect 25161 1074 25167 1108
rect 25121 1036 25167 1074
rect 25121 1002 25127 1036
rect 25161 1002 25167 1036
rect 25121 990 25167 1002
rect 25251 1108 25297 1113
rect 25251 1074 25257 1108
rect 25291 1074 25297 1108
rect 25251 1036 25297 1074
rect 25251 1002 25257 1036
rect 25291 1002 25297 1036
rect 25251 990 25297 1002
rect 25381 1108 25427 1146
rect 25497 1189 25571 1213
rect 25497 1137 25508 1189
rect 25560 1137 25571 1189
rect 25497 1113 25571 1137
rect 25627 1189 25701 1213
rect 25627 1137 25638 1189
rect 25690 1137 25701 1189
rect 25627 1113 25701 1137
rect 25771 1180 25817 1218
rect 25901 1324 25947 1336
rect 25901 1290 25907 1324
rect 25941 1290 25947 1324
rect 25901 1252 25947 1290
rect 25901 1218 25907 1252
rect 25941 1218 25947 1252
rect 25901 1213 25947 1218
rect 26031 1324 26077 1336
rect 26031 1290 26037 1324
rect 26071 1290 26077 1324
rect 26031 1252 26077 1290
rect 26031 1218 26037 1252
rect 26071 1218 26077 1252
rect 26031 1213 26077 1218
rect 26161 1324 26207 1550
rect 26412 1872 26476 1884
rect 26412 1865 26427 1872
rect 26461 1865 26476 1872
rect 26412 1813 26418 1865
rect 26470 1813 26476 1865
rect 26412 1801 26476 1813
rect 26412 1749 26418 1801
rect 26470 1749 26476 1801
rect 26412 1737 26476 1749
rect 26412 1685 26418 1737
rect 26470 1685 26476 1737
rect 26412 1673 26476 1685
rect 26412 1621 26418 1673
rect 26470 1621 26476 1673
rect 26412 1609 26476 1621
rect 26412 1557 26418 1609
rect 26470 1557 26476 1609
rect 26412 1550 26427 1557
rect 26461 1550 26476 1557
rect 26412 1538 26476 1550
rect 26551 1872 26597 1884
rect 26551 1838 26557 1872
rect 26591 1838 26597 1872
rect 26551 1800 26597 1838
rect 26551 1766 26557 1800
rect 26591 1766 26597 1800
rect 26551 1728 26597 1766
rect 26551 1694 26557 1728
rect 26591 1694 26597 1728
rect 26551 1656 26597 1694
rect 26551 1622 26557 1656
rect 26591 1622 26597 1656
rect 26551 1584 26597 1622
rect 26551 1550 26557 1584
rect 26591 1550 26597 1584
rect 26161 1290 26167 1324
rect 26201 1290 26207 1324
rect 26161 1252 26207 1290
rect 26161 1218 26167 1252
rect 26201 1218 26207 1252
rect 25771 1146 25777 1180
rect 25811 1146 25817 1180
rect 25381 1074 25387 1108
rect 25421 1074 25427 1108
rect 25381 1036 25427 1074
rect 25381 1002 25387 1036
rect 25421 1002 25427 1036
rect 25381 990 25427 1002
rect 25511 1108 25557 1113
rect 25511 1074 25517 1108
rect 25551 1074 25557 1108
rect 25511 1036 25557 1074
rect 25511 1002 25517 1036
rect 25551 1002 25557 1036
rect 25511 990 25557 1002
rect 25641 1108 25687 1113
rect 25641 1074 25647 1108
rect 25681 1074 25687 1108
rect 25641 1036 25687 1074
rect 25641 1002 25647 1036
rect 25681 1002 25687 1036
rect 25641 990 25687 1002
rect 25771 1108 25817 1146
rect 25887 1189 25961 1213
rect 25887 1137 25898 1189
rect 25950 1137 25961 1189
rect 25887 1113 25961 1137
rect 26017 1189 26091 1213
rect 26017 1137 26028 1189
rect 26080 1137 26091 1189
rect 26017 1113 26091 1137
rect 26161 1180 26207 1218
rect 26291 1324 26337 1336
rect 26291 1290 26297 1324
rect 26331 1290 26337 1324
rect 26291 1252 26337 1290
rect 26291 1218 26297 1252
rect 26331 1218 26337 1252
rect 26291 1213 26337 1218
rect 26421 1324 26467 1336
rect 26421 1290 26427 1324
rect 26461 1290 26467 1324
rect 26421 1252 26467 1290
rect 26421 1218 26427 1252
rect 26461 1218 26467 1252
rect 26421 1213 26467 1218
rect 26551 1324 26597 1550
rect 26802 1872 26866 1884
rect 26802 1865 26817 1872
rect 26851 1865 26866 1872
rect 26802 1813 26808 1865
rect 26860 1813 26866 1865
rect 26802 1801 26866 1813
rect 26802 1749 26808 1801
rect 26860 1749 26866 1801
rect 26802 1737 26866 1749
rect 26802 1685 26808 1737
rect 26860 1685 26866 1737
rect 26802 1673 26866 1685
rect 26802 1621 26808 1673
rect 26860 1621 26866 1673
rect 26802 1609 26866 1621
rect 26802 1557 26808 1609
rect 26860 1557 26866 1609
rect 26802 1550 26817 1557
rect 26851 1550 26866 1557
rect 26802 1538 26866 1550
rect 26941 1872 26987 1884
rect 26941 1838 26947 1872
rect 26981 1838 26987 1872
rect 26941 1800 26987 1838
rect 26941 1766 26947 1800
rect 26981 1766 26987 1800
rect 26941 1728 26987 1766
rect 26941 1694 26947 1728
rect 26981 1694 26987 1728
rect 26941 1656 26987 1694
rect 26941 1622 26947 1656
rect 26981 1622 26987 1656
rect 26941 1584 26987 1622
rect 26941 1550 26947 1584
rect 26981 1550 26987 1584
rect 26551 1290 26557 1324
rect 26591 1290 26597 1324
rect 26551 1252 26597 1290
rect 26551 1218 26557 1252
rect 26591 1218 26597 1252
rect 26161 1146 26167 1180
rect 26201 1146 26207 1180
rect 25771 1074 25777 1108
rect 25811 1074 25817 1108
rect 25771 1036 25817 1074
rect 25771 1002 25777 1036
rect 25811 1002 25817 1036
rect 25771 990 25817 1002
rect 25901 1108 25947 1113
rect 25901 1074 25907 1108
rect 25941 1074 25947 1108
rect 25901 1036 25947 1074
rect 25901 1002 25907 1036
rect 25941 1002 25947 1036
rect 25901 990 25947 1002
rect 26031 1108 26077 1113
rect 26031 1074 26037 1108
rect 26071 1074 26077 1108
rect 26031 1036 26077 1074
rect 26031 1002 26037 1036
rect 26071 1002 26077 1036
rect 26031 990 26077 1002
rect 26161 1108 26207 1146
rect 26277 1189 26351 1213
rect 26277 1137 26288 1189
rect 26340 1137 26351 1189
rect 26277 1113 26351 1137
rect 26407 1189 26481 1213
rect 26407 1137 26418 1189
rect 26470 1137 26481 1189
rect 26407 1113 26481 1137
rect 26551 1180 26597 1218
rect 26681 1324 26727 1336
rect 26681 1290 26687 1324
rect 26721 1290 26727 1324
rect 26681 1252 26727 1290
rect 26681 1218 26687 1252
rect 26721 1218 26727 1252
rect 26681 1213 26727 1218
rect 26811 1324 26857 1336
rect 26811 1290 26817 1324
rect 26851 1290 26857 1324
rect 26811 1252 26857 1290
rect 26811 1218 26817 1252
rect 26851 1218 26857 1252
rect 26811 1213 26857 1218
rect 26941 1324 26987 1550
rect 26941 1290 26947 1324
rect 26981 1290 26987 1324
rect 26941 1252 26987 1290
rect 26941 1218 26947 1252
rect 26981 1218 26987 1252
rect 26551 1146 26557 1180
rect 26591 1146 26597 1180
rect 26161 1074 26167 1108
rect 26201 1074 26207 1108
rect 26161 1036 26207 1074
rect 26161 1002 26167 1036
rect 26201 1002 26207 1036
rect 26161 990 26207 1002
rect 26291 1108 26337 1113
rect 26291 1074 26297 1108
rect 26331 1074 26337 1108
rect 26291 1036 26337 1074
rect 26291 1002 26297 1036
rect 26331 1002 26337 1036
rect 26291 990 26337 1002
rect 26421 1108 26467 1113
rect 26421 1074 26427 1108
rect 26461 1074 26467 1108
rect 26421 1036 26467 1074
rect 26421 1002 26427 1036
rect 26461 1002 26467 1036
rect 26421 990 26467 1002
rect 26551 1108 26597 1146
rect 26667 1189 26741 1213
rect 26667 1137 26678 1189
rect 26730 1137 26741 1189
rect 26667 1113 26741 1137
rect 26797 1189 26871 1213
rect 26797 1137 26808 1189
rect 26860 1137 26871 1189
rect 26797 1113 26871 1137
rect 26941 1180 26987 1218
rect 27071 1324 27117 1336
rect 27071 1290 27077 1324
rect 27111 1290 27117 1324
rect 27071 1252 27117 1290
rect 27071 1218 27077 1252
rect 27111 1218 27117 1252
rect 27071 1213 27117 1218
rect 26941 1146 26947 1180
rect 26981 1146 26987 1180
rect 26551 1074 26557 1108
rect 26591 1074 26597 1108
rect 26551 1036 26597 1074
rect 26551 1002 26557 1036
rect 26591 1002 26597 1036
rect 26551 990 26597 1002
rect 26681 1108 26727 1113
rect 26681 1074 26687 1108
rect 26721 1074 26727 1108
rect 26681 1036 26727 1074
rect 26681 1002 26687 1036
rect 26721 1002 26727 1036
rect 26681 990 26727 1002
rect 26811 1108 26857 1113
rect 26811 1074 26817 1108
rect 26851 1074 26857 1108
rect 26811 1036 26857 1074
rect 26811 1002 26817 1036
rect 26851 1002 26857 1036
rect 26811 990 26857 1002
rect 26941 1108 26987 1146
rect 27057 1189 27131 1213
rect 27057 1137 27068 1189
rect 27120 1137 27131 1189
rect 27057 1113 27131 1137
rect 26941 1074 26947 1108
rect 26981 1074 26987 1108
rect 26941 1036 26987 1074
rect 26941 1002 26947 1036
rect 26981 1002 26987 1036
rect 26941 990 26987 1002
rect 27071 1108 27117 1113
rect 27071 1074 27077 1108
rect 27111 1074 27117 1108
rect 27071 1036 27117 1074
rect 27071 1002 27077 1036
rect 27111 1002 27117 1036
rect 27071 990 27117 1002
rect 12493 916 12567 923
rect 12493 864 12504 916
rect 12556 864 12567 916
rect 13320 916 13394 923
rect 12493 857 12567 864
rect 13190 907 13264 913
rect 13190 873 13210 907
rect 13244 873 13264 907
rect 13190 797 13264 873
rect 13320 864 13331 916
rect 13383 864 13394 916
rect 13710 916 13784 923
rect 13320 857 13394 864
rect 13450 907 13524 913
rect 13450 873 13470 907
rect 13504 873 13524 907
rect 13450 797 13524 873
rect 13580 907 13654 913
rect 13580 873 13600 907
rect 13634 873 13654 907
rect 13580 797 13654 873
rect 13710 864 13721 916
rect 13773 864 13784 916
rect 14100 916 14174 923
rect 13710 857 13784 864
rect 13840 907 13914 913
rect 13840 873 13860 907
rect 13894 873 13914 907
rect 13840 797 13914 873
rect 13970 907 14044 913
rect 13970 873 13990 907
rect 14024 873 14044 907
rect 13970 797 14044 873
rect 14100 864 14111 916
rect 14163 864 14174 916
rect 14490 916 14564 923
rect 14100 857 14174 864
rect 14230 907 14304 913
rect 14230 873 14250 907
rect 14284 873 14304 907
rect 14230 797 14304 873
rect 14360 907 14434 913
rect 14360 873 14380 907
rect 14414 873 14434 907
rect 14360 797 14434 873
rect 14490 864 14501 916
rect 14553 864 14564 916
rect 14880 916 14954 923
rect 14490 857 14564 864
rect 14620 907 14694 913
rect 14620 873 14640 907
rect 14674 873 14694 907
rect 14620 797 14694 873
rect 14750 907 14824 913
rect 14750 873 14770 907
rect 14804 873 14824 907
rect 14750 797 14824 873
rect 14880 864 14891 916
rect 14943 864 14954 916
rect 15270 916 15344 923
rect 14880 857 14954 864
rect 15010 907 15084 913
rect 15010 873 15030 907
rect 15064 873 15084 907
rect 15010 797 15084 873
rect 15140 907 15214 913
rect 15140 873 15160 907
rect 15194 873 15214 907
rect 15140 797 15214 873
rect 15270 864 15281 916
rect 15333 864 15344 916
rect 24085 916 24159 923
rect 15270 857 15344 864
rect 15400 907 15474 913
rect 15400 873 15420 907
rect 15454 873 15474 907
rect 15400 797 15474 873
rect 24085 864 24096 916
rect 24148 864 24159 916
rect 24912 916 24986 923
rect 24085 857 24159 864
rect 24782 907 24856 913
rect 24782 873 24802 907
rect 24836 873 24856 907
rect 24782 797 24856 873
rect 24912 864 24923 916
rect 24975 864 24986 916
rect 25302 916 25376 923
rect 24912 857 24986 864
rect 25042 907 25116 913
rect 25042 873 25062 907
rect 25096 873 25116 907
rect 25042 797 25116 873
rect 25172 907 25246 913
rect 25172 873 25192 907
rect 25226 873 25246 907
rect 25172 797 25246 873
rect 25302 864 25313 916
rect 25365 864 25376 916
rect 25692 916 25766 923
rect 25302 857 25376 864
rect 25432 907 25506 913
rect 25432 873 25452 907
rect 25486 873 25506 907
rect 25432 797 25506 873
rect 25562 907 25636 913
rect 25562 873 25582 907
rect 25616 873 25636 907
rect 25562 797 25636 873
rect 25692 864 25703 916
rect 25755 864 25766 916
rect 26082 916 26156 923
rect 25692 857 25766 864
rect 25822 907 25896 913
rect 25822 873 25842 907
rect 25876 873 25896 907
rect 25822 797 25896 873
rect 25952 907 26026 913
rect 25952 873 25972 907
rect 26006 873 26026 907
rect 25952 797 26026 873
rect 26082 864 26093 916
rect 26145 864 26156 916
rect 26472 916 26546 923
rect 26082 857 26156 864
rect 26212 907 26286 913
rect 26212 873 26232 907
rect 26266 873 26286 907
rect 26212 797 26286 873
rect 26342 907 26416 913
rect 26342 873 26362 907
rect 26396 873 26416 907
rect 26342 797 26416 873
rect 26472 864 26483 916
rect 26535 864 26546 916
rect 26862 916 26936 923
rect 26472 857 26546 864
rect 26602 907 26676 913
rect 26602 873 26622 907
rect 26656 873 26676 907
rect 26602 797 26676 873
rect 26732 907 26806 913
rect 26732 873 26752 907
rect 26786 873 26806 907
rect 26732 797 26806 873
rect 26862 864 26873 916
rect 26925 864 26936 916
rect 26862 857 26936 864
rect 26992 907 27066 913
rect 26992 873 27012 907
rect 27046 873 27066 907
rect 26992 797 27066 873
rect 12823 783 15697 797
rect 12823 731 12833 783
rect 12885 731 12897 783
rect 12949 731 12961 783
rect 13013 774 13657 783
rect 13013 740 13196 774
rect 13230 740 13268 774
rect 13302 740 13340 774
rect 13374 740 13412 774
rect 13446 740 13484 774
rect 13518 740 13586 774
rect 13620 740 13657 774
rect 13013 731 13657 740
rect 13709 731 13721 783
rect 13773 731 13785 783
rect 13837 774 14437 783
rect 13837 740 13874 774
rect 13908 740 13976 774
rect 14010 740 14048 774
rect 14082 740 14120 774
rect 14154 740 14192 774
rect 14226 740 14264 774
rect 14298 740 14366 774
rect 14400 740 14437 774
rect 13837 731 14437 740
rect 14489 731 14501 783
rect 14553 731 14565 783
rect 14617 774 15217 783
rect 14617 740 14654 774
rect 14688 740 14756 774
rect 14790 740 14828 774
rect 14862 740 14900 774
rect 14934 740 14972 774
rect 15006 740 15044 774
rect 15078 740 15146 774
rect 15180 740 15217 774
rect 14617 731 15217 740
rect 15269 731 15281 783
rect 15333 731 15345 783
rect 15397 774 15697 783
rect 15397 740 15434 774
rect 15468 740 15697 774
rect 15397 731 15697 740
rect 12823 717 15697 731
rect 24415 783 27289 797
rect 24415 731 24425 783
rect 24477 731 24489 783
rect 24541 731 24553 783
rect 24605 774 25249 783
rect 24605 740 24788 774
rect 24822 740 24860 774
rect 24894 740 24932 774
rect 24966 740 25004 774
rect 25038 740 25076 774
rect 25110 740 25178 774
rect 25212 740 25249 774
rect 24605 731 25249 740
rect 25301 731 25313 783
rect 25365 731 25377 783
rect 25429 774 26029 783
rect 25429 740 25466 774
rect 25500 740 25568 774
rect 25602 740 25640 774
rect 25674 740 25712 774
rect 25746 740 25784 774
rect 25818 740 25856 774
rect 25890 740 25958 774
rect 25992 740 26029 774
rect 25429 731 26029 740
rect 26081 731 26093 783
rect 26145 731 26157 783
rect 26209 774 26809 783
rect 26209 740 26246 774
rect 26280 740 26348 774
rect 26382 740 26420 774
rect 26454 740 26492 774
rect 26526 740 26564 774
rect 26598 740 26636 774
rect 26670 740 26738 774
rect 26772 740 26809 774
rect 26209 731 26809 740
rect 26861 731 26873 783
rect 26925 731 26937 783
rect 26989 774 27289 783
rect 26989 740 27026 774
rect 27060 740 27289 774
rect 26989 731 27289 740
rect 24415 717 27289 731
<< via1 >>
rect 12833 5443 12885 5495
rect 12897 5443 12949 5495
rect 12961 5443 13013 5495
rect 13657 5486 13709 5495
rect 13657 5452 13658 5486
rect 13658 5452 13692 5486
rect 13692 5452 13709 5486
rect 13657 5443 13709 5452
rect 13721 5486 13773 5495
rect 13721 5452 13730 5486
rect 13730 5452 13764 5486
rect 13764 5452 13773 5486
rect 13721 5443 13773 5452
rect 13785 5486 13837 5495
rect 14437 5486 14489 5495
rect 13785 5452 13802 5486
rect 13802 5452 13836 5486
rect 13836 5452 13837 5486
rect 14437 5452 14438 5486
rect 14438 5452 14472 5486
rect 14472 5452 14489 5486
rect 13785 5443 13837 5452
rect 14437 5443 14489 5452
rect 14501 5486 14553 5495
rect 14501 5452 14510 5486
rect 14510 5452 14544 5486
rect 14544 5452 14553 5486
rect 14501 5443 14553 5452
rect 14565 5486 14617 5495
rect 14565 5452 14582 5486
rect 14582 5452 14616 5486
rect 14616 5452 14617 5486
rect 14565 5443 14617 5452
rect 15217 5443 15269 5495
rect 15281 5443 15333 5495
rect 15345 5443 15397 5495
rect 24425 5443 24477 5495
rect 24489 5443 24541 5495
rect 24553 5443 24605 5495
rect 25249 5486 25301 5495
rect 25249 5452 25250 5486
rect 25250 5452 25284 5486
rect 25284 5452 25301 5486
rect 25249 5443 25301 5452
rect 25313 5486 25365 5495
rect 25313 5452 25322 5486
rect 25322 5452 25356 5486
rect 25356 5452 25365 5486
rect 25313 5443 25365 5452
rect 25377 5486 25429 5495
rect 26029 5486 26081 5495
rect 25377 5452 25394 5486
rect 25394 5452 25428 5486
rect 25428 5452 25429 5486
rect 26029 5452 26030 5486
rect 26030 5452 26064 5486
rect 26064 5452 26081 5486
rect 25377 5443 25429 5452
rect 26029 5443 26081 5452
rect 26093 5486 26145 5495
rect 26093 5452 26102 5486
rect 26102 5452 26136 5486
rect 26136 5452 26145 5486
rect 26093 5443 26145 5452
rect 26157 5486 26209 5495
rect 26157 5452 26174 5486
rect 26174 5452 26208 5486
rect 26208 5452 26209 5486
rect 26157 5443 26209 5452
rect 26809 5443 26861 5495
rect 26873 5443 26925 5495
rect 26937 5443 26989 5495
rect 12504 5310 12556 5362
rect 13009 5310 13061 5362
rect 13073 5353 13125 5362
rect 13073 5319 13080 5353
rect 13080 5319 13114 5353
rect 13114 5319 13125 5353
rect 13073 5310 13125 5319
rect 13331 5353 13383 5362
rect 13331 5319 13340 5353
rect 13340 5319 13374 5353
rect 13374 5319 13383 5353
rect 13331 5310 13383 5319
rect 13721 5353 13773 5362
rect 13721 5319 13730 5353
rect 13730 5319 13764 5353
rect 13764 5319 13773 5353
rect 13721 5310 13773 5319
rect 14111 5353 14163 5362
rect 14111 5319 14120 5353
rect 14120 5319 14154 5353
rect 14154 5319 14163 5353
rect 14111 5310 14163 5319
rect 14501 5353 14553 5362
rect 14501 5319 14510 5353
rect 14510 5319 14544 5353
rect 14544 5319 14553 5353
rect 14501 5310 14553 5319
rect 14891 5353 14943 5362
rect 14891 5319 14900 5353
rect 14900 5319 14934 5353
rect 14934 5319 14943 5353
rect 14891 5310 14943 5319
rect 24096 5310 24148 5362
rect 24601 5310 24653 5362
rect 24665 5353 24717 5362
rect 24665 5319 24672 5353
rect 24672 5319 24706 5353
rect 24706 5319 24717 5353
rect 24665 5310 24717 5319
rect 24923 5353 24975 5362
rect 24923 5319 24932 5353
rect 24932 5319 24966 5353
rect 24966 5319 24975 5353
rect 24923 5310 24975 5319
rect 25313 5353 25365 5362
rect 25313 5319 25322 5353
rect 25322 5319 25356 5353
rect 25356 5319 25365 5353
rect 25313 5310 25365 5319
rect 25703 5353 25755 5362
rect 25703 5319 25712 5353
rect 25712 5319 25746 5353
rect 25746 5319 25755 5353
rect 25703 5310 25755 5319
rect 26093 5353 26145 5362
rect 26093 5319 26102 5353
rect 26102 5319 26136 5353
rect 26136 5319 26145 5353
rect 26093 5310 26145 5319
rect 26483 5353 26535 5362
rect 26483 5319 26492 5353
rect 26492 5319 26526 5353
rect 26526 5319 26535 5353
rect 26483 5310 26535 5319
rect 13006 5190 13015 5217
rect 13015 5190 13049 5217
rect 13049 5190 13058 5217
rect 13006 5165 13058 5190
rect 13006 5152 13058 5153
rect 13006 5118 13015 5152
rect 13015 5118 13049 5152
rect 13049 5118 13058 5152
rect 13006 5101 13058 5118
rect 13006 5080 13058 5089
rect 13006 5046 13015 5080
rect 13015 5046 13049 5080
rect 13049 5046 13058 5080
rect 13006 5037 13058 5046
rect 13006 5008 13058 5025
rect 13006 4974 13015 5008
rect 13015 4974 13049 5008
rect 13049 4974 13058 5008
rect 13006 4973 13058 4974
rect 13136 5080 13188 5089
rect 13136 5046 13145 5080
rect 13145 5046 13179 5080
rect 13179 5046 13188 5080
rect 13136 5037 13188 5046
rect 13006 4936 13058 4961
rect 13006 4909 13015 4936
rect 13015 4909 13049 4936
rect 13049 4909 13058 4936
rect 13396 5080 13448 5089
rect 13396 5046 13405 5080
rect 13405 5046 13439 5080
rect 13439 5046 13448 5080
rect 13396 5037 13448 5046
rect 13526 5080 13578 5089
rect 13526 5046 13535 5080
rect 13535 5046 13569 5080
rect 13569 5046 13578 5080
rect 13526 5037 13578 5046
rect 13786 5080 13838 5089
rect 13786 5046 13795 5080
rect 13795 5046 13829 5080
rect 13829 5046 13838 5080
rect 13786 5037 13838 5046
rect 13916 5080 13968 5089
rect 13916 5046 13925 5080
rect 13925 5046 13959 5080
rect 13959 5046 13968 5080
rect 13916 5037 13968 5046
rect 13396 4642 13405 4669
rect 13405 4642 13439 4669
rect 13439 4642 13448 4669
rect 13396 4617 13448 4642
rect 13396 4604 13448 4605
rect 13396 4570 13405 4604
rect 13405 4570 13439 4604
rect 13439 4570 13448 4604
rect 13396 4553 13448 4570
rect 13396 4532 13448 4541
rect 13396 4498 13405 4532
rect 13405 4498 13439 4532
rect 13439 4498 13448 4532
rect 13396 4489 13448 4498
rect 13396 4460 13448 4477
rect 13396 4426 13405 4460
rect 13405 4426 13439 4460
rect 13439 4426 13448 4460
rect 13396 4425 13448 4426
rect 13396 4388 13448 4413
rect 13396 4361 13405 4388
rect 13405 4361 13439 4388
rect 13439 4361 13448 4388
rect 14176 5080 14228 5089
rect 14176 5046 14185 5080
rect 14185 5046 14219 5080
rect 14219 5046 14228 5080
rect 14176 5037 14228 5046
rect 14306 5080 14358 5089
rect 14306 5046 14315 5080
rect 14315 5046 14349 5080
rect 14349 5046 14358 5080
rect 14306 5037 14358 5046
rect 13786 4642 13795 4669
rect 13795 4642 13829 4669
rect 13829 4642 13838 4669
rect 13786 4617 13838 4642
rect 13786 4604 13838 4605
rect 13786 4570 13795 4604
rect 13795 4570 13829 4604
rect 13829 4570 13838 4604
rect 13786 4553 13838 4570
rect 13786 4532 13838 4541
rect 13786 4498 13795 4532
rect 13795 4498 13829 4532
rect 13829 4498 13838 4532
rect 13786 4489 13838 4498
rect 13786 4460 13838 4477
rect 13786 4426 13795 4460
rect 13795 4426 13829 4460
rect 13829 4426 13838 4460
rect 13786 4425 13838 4426
rect 13786 4388 13838 4413
rect 13786 4361 13795 4388
rect 13795 4361 13829 4388
rect 13829 4361 13838 4388
rect 14566 5080 14618 5089
rect 14566 5046 14575 5080
rect 14575 5046 14609 5080
rect 14609 5046 14618 5080
rect 14566 5037 14618 5046
rect 14696 5080 14748 5089
rect 14696 5046 14705 5080
rect 14705 5046 14739 5080
rect 14739 5046 14748 5080
rect 14696 5037 14748 5046
rect 24598 5190 24607 5217
rect 24607 5190 24641 5217
rect 24641 5190 24650 5217
rect 24598 5165 24650 5190
rect 14176 4642 14185 4669
rect 14185 4642 14219 4669
rect 14219 4642 14228 4669
rect 14176 4617 14228 4642
rect 14176 4604 14228 4605
rect 14176 4570 14185 4604
rect 14185 4570 14219 4604
rect 14219 4570 14228 4604
rect 14176 4553 14228 4570
rect 14176 4532 14228 4541
rect 14176 4498 14185 4532
rect 14185 4498 14219 4532
rect 14219 4498 14228 4532
rect 14176 4489 14228 4498
rect 14176 4460 14228 4477
rect 14176 4426 14185 4460
rect 14185 4426 14219 4460
rect 14219 4426 14228 4460
rect 14176 4425 14228 4426
rect 14176 4388 14228 4413
rect 14176 4361 14185 4388
rect 14185 4361 14219 4388
rect 14219 4361 14228 4388
rect 14956 5080 15008 5089
rect 14956 5046 14965 5080
rect 14965 5046 14999 5080
rect 14999 5046 15008 5080
rect 14956 5037 15008 5046
rect 15086 5080 15138 5089
rect 15086 5046 15095 5080
rect 15095 5046 15129 5080
rect 15129 5046 15138 5080
rect 15086 5037 15138 5046
rect 24598 5152 24650 5153
rect 24598 5118 24607 5152
rect 24607 5118 24641 5152
rect 24641 5118 24650 5152
rect 24598 5101 24650 5118
rect 24598 5080 24650 5089
rect 24598 5046 24607 5080
rect 24607 5046 24641 5080
rect 24641 5046 24650 5080
rect 24598 5037 24650 5046
rect 14566 4642 14575 4669
rect 14575 4642 14609 4669
rect 14609 4642 14618 4669
rect 14566 4617 14618 4642
rect 14566 4604 14618 4605
rect 14566 4570 14575 4604
rect 14575 4570 14609 4604
rect 14609 4570 14618 4604
rect 14566 4553 14618 4570
rect 14566 4532 14618 4541
rect 14566 4498 14575 4532
rect 14575 4498 14609 4532
rect 14609 4498 14618 4532
rect 14566 4489 14618 4498
rect 14566 4460 14618 4477
rect 14566 4426 14575 4460
rect 14575 4426 14609 4460
rect 14609 4426 14618 4460
rect 14566 4425 14618 4426
rect 14566 4388 14618 4413
rect 14566 4361 14575 4388
rect 14575 4361 14609 4388
rect 14609 4361 14618 4388
rect 24598 5008 24650 5025
rect 24598 4974 24607 5008
rect 24607 4974 24641 5008
rect 24641 4974 24650 5008
rect 24598 4973 24650 4974
rect 24728 5080 24780 5089
rect 24728 5046 24737 5080
rect 24737 5046 24771 5080
rect 24771 5046 24780 5080
rect 24728 5037 24780 5046
rect 15317 4915 15369 4924
rect 15317 4881 15349 4915
rect 15349 4881 15369 4915
rect 15317 4872 15369 4881
rect 15381 4915 15433 4924
rect 15381 4881 15387 4915
rect 15387 4881 15421 4915
rect 15421 4881 15433 4915
rect 15381 4872 15433 4881
rect 15445 4915 15497 4924
rect 15445 4881 15459 4915
rect 15459 4881 15493 4915
rect 15493 4881 15497 4915
rect 15445 4872 15497 4881
rect 24598 4936 24650 4961
rect 24598 4909 24607 4936
rect 24607 4909 24641 4936
rect 24641 4909 24650 4936
rect 24988 5080 25040 5089
rect 24988 5046 24997 5080
rect 24997 5046 25031 5080
rect 25031 5046 25040 5080
rect 24988 5037 25040 5046
rect 25118 5080 25170 5089
rect 25118 5046 25127 5080
rect 25127 5046 25161 5080
rect 25161 5046 25170 5080
rect 25118 5037 25170 5046
rect 15204 4781 15256 4833
rect 14956 4642 14965 4669
rect 14965 4642 14999 4669
rect 14999 4642 15008 4669
rect 14956 4617 15008 4642
rect 14956 4604 15008 4605
rect 14956 4570 14965 4604
rect 14965 4570 14999 4604
rect 14999 4570 15008 4604
rect 14956 4553 15008 4570
rect 14956 4532 15008 4541
rect 14956 4498 14965 4532
rect 14965 4498 14999 4532
rect 14999 4498 15008 4532
rect 14956 4489 15008 4498
rect 14956 4460 15008 4477
rect 14956 4426 14965 4460
rect 14965 4426 14999 4460
rect 14999 4426 15008 4460
rect 14956 4425 15008 4426
rect 14956 4388 15008 4413
rect 14956 4361 14965 4388
rect 14965 4361 14999 4388
rect 14999 4361 15008 4388
rect 15290 4676 15342 4685
rect 15290 4642 15299 4676
rect 15299 4642 15333 4676
rect 15333 4642 15342 4676
rect 15290 4633 15342 4642
rect 15200 4388 15252 4397
rect 15200 4354 15209 4388
rect 15209 4354 15243 4388
rect 15243 4354 15252 4388
rect 15200 4345 15252 4354
rect 15470 4676 15522 4685
rect 15470 4642 15479 4676
rect 15479 4642 15513 4676
rect 15513 4642 15522 4676
rect 15470 4633 15522 4642
rect 15380 4388 15432 4391
rect 15380 4354 15389 4388
rect 15389 4354 15423 4388
rect 15423 4354 15432 4388
rect 15380 4339 15432 4354
rect 25378 5080 25430 5089
rect 25378 5046 25387 5080
rect 25387 5046 25421 5080
rect 25421 5046 25430 5080
rect 25378 5037 25430 5046
rect 25508 5080 25560 5089
rect 25508 5046 25517 5080
rect 25517 5046 25551 5080
rect 25551 5046 25560 5080
rect 25508 5037 25560 5046
rect 15560 4388 15612 4391
rect 15560 4354 15569 4388
rect 15569 4354 15603 4388
rect 15603 4354 15612 4388
rect 15560 4339 15612 4354
rect 24988 4642 24997 4669
rect 24997 4642 25031 4669
rect 25031 4642 25040 4669
rect 24988 4617 25040 4642
rect 24988 4604 25040 4605
rect 24988 4570 24997 4604
rect 24997 4570 25031 4604
rect 25031 4570 25040 4604
rect 24988 4553 25040 4570
rect 24988 4532 25040 4541
rect 24988 4498 24997 4532
rect 24997 4498 25031 4532
rect 25031 4498 25040 4532
rect 24988 4489 25040 4498
rect 24988 4460 25040 4477
rect 24988 4426 24997 4460
rect 24997 4426 25031 4460
rect 25031 4426 25040 4460
rect 24988 4425 25040 4426
rect 24988 4388 25040 4413
rect 24988 4361 24997 4388
rect 24997 4361 25031 4388
rect 25031 4361 25040 4388
rect 25768 5080 25820 5089
rect 25768 5046 25777 5080
rect 25777 5046 25811 5080
rect 25811 5046 25820 5080
rect 25768 5037 25820 5046
rect 25898 5080 25950 5089
rect 25898 5046 25907 5080
rect 25907 5046 25941 5080
rect 25941 5046 25950 5080
rect 25898 5037 25950 5046
rect 25378 4642 25387 4669
rect 25387 4642 25421 4669
rect 25421 4642 25430 4669
rect 25378 4617 25430 4642
rect 25378 4604 25430 4605
rect 25378 4570 25387 4604
rect 25387 4570 25421 4604
rect 25421 4570 25430 4604
rect 25378 4553 25430 4570
rect 25378 4532 25430 4541
rect 25378 4498 25387 4532
rect 25387 4498 25421 4532
rect 25421 4498 25430 4532
rect 25378 4489 25430 4498
rect 25378 4460 25430 4477
rect 25378 4426 25387 4460
rect 25387 4426 25421 4460
rect 25421 4426 25430 4460
rect 25378 4425 25430 4426
rect 25378 4388 25430 4413
rect 25378 4361 25387 4388
rect 25387 4361 25421 4388
rect 25421 4361 25430 4388
rect 26158 5080 26210 5089
rect 26158 5046 26167 5080
rect 26167 5046 26201 5080
rect 26201 5046 26210 5080
rect 26158 5037 26210 5046
rect 26288 5080 26340 5089
rect 26288 5046 26297 5080
rect 26297 5046 26331 5080
rect 26331 5046 26340 5080
rect 26288 5037 26340 5046
rect 25768 4642 25777 4669
rect 25777 4642 25811 4669
rect 25811 4642 25820 4669
rect 25768 4617 25820 4642
rect 25768 4604 25820 4605
rect 25768 4570 25777 4604
rect 25777 4570 25811 4604
rect 25811 4570 25820 4604
rect 25768 4553 25820 4570
rect 25768 4532 25820 4541
rect 25768 4498 25777 4532
rect 25777 4498 25811 4532
rect 25811 4498 25820 4532
rect 25768 4489 25820 4498
rect 25768 4460 25820 4477
rect 25768 4426 25777 4460
rect 25777 4426 25811 4460
rect 25811 4426 25820 4460
rect 25768 4425 25820 4426
rect 25768 4388 25820 4413
rect 25768 4361 25777 4388
rect 25777 4361 25811 4388
rect 25811 4361 25820 4388
rect 26548 5080 26600 5089
rect 26548 5046 26557 5080
rect 26557 5046 26591 5080
rect 26591 5046 26600 5080
rect 26548 5037 26600 5046
rect 26678 5080 26730 5089
rect 26678 5046 26687 5080
rect 26687 5046 26721 5080
rect 26721 5046 26730 5080
rect 26678 5037 26730 5046
rect 26158 4642 26167 4669
rect 26167 4642 26201 4669
rect 26201 4642 26210 4669
rect 26158 4617 26210 4642
rect 26158 4604 26210 4605
rect 26158 4570 26167 4604
rect 26167 4570 26201 4604
rect 26201 4570 26210 4604
rect 26158 4553 26210 4570
rect 26158 4532 26210 4541
rect 26158 4498 26167 4532
rect 26167 4498 26201 4532
rect 26201 4498 26210 4532
rect 26158 4489 26210 4498
rect 26158 4460 26210 4477
rect 26158 4426 26167 4460
rect 26167 4426 26201 4460
rect 26201 4426 26210 4460
rect 26158 4425 26210 4426
rect 26158 4388 26210 4413
rect 26158 4361 26167 4388
rect 26167 4361 26201 4388
rect 26201 4361 26210 4388
rect 26909 4915 26961 4924
rect 26909 4881 26941 4915
rect 26941 4881 26961 4915
rect 26909 4872 26961 4881
rect 26973 4915 27025 4924
rect 26973 4881 26979 4915
rect 26979 4881 27013 4915
rect 27013 4881 27025 4915
rect 26973 4872 27025 4881
rect 27037 4915 27089 4924
rect 27037 4881 27051 4915
rect 27051 4881 27085 4915
rect 27085 4881 27089 4915
rect 27037 4872 27089 4881
rect 26796 4781 26848 4833
rect 26548 4642 26557 4669
rect 26557 4642 26591 4669
rect 26591 4642 26600 4669
rect 26548 4617 26600 4642
rect 26548 4604 26600 4605
rect 26548 4570 26557 4604
rect 26557 4570 26591 4604
rect 26591 4570 26600 4604
rect 26548 4553 26600 4570
rect 26548 4532 26600 4541
rect 26548 4498 26557 4532
rect 26557 4498 26591 4532
rect 26591 4498 26600 4532
rect 26548 4489 26600 4498
rect 26548 4460 26600 4477
rect 26548 4426 26557 4460
rect 26557 4426 26591 4460
rect 26591 4426 26600 4460
rect 26548 4425 26600 4426
rect 26548 4388 26600 4413
rect 26548 4361 26557 4388
rect 26557 4361 26591 4388
rect 26591 4361 26600 4388
rect 26882 4676 26934 4685
rect 26882 4642 26891 4676
rect 26891 4642 26925 4676
rect 26925 4642 26934 4676
rect 26882 4633 26934 4642
rect 26792 4388 26844 4397
rect 26792 4354 26801 4388
rect 26801 4354 26835 4388
rect 26835 4354 26844 4388
rect 26792 4345 26844 4354
rect 27062 4676 27114 4685
rect 27062 4642 27071 4676
rect 27071 4642 27105 4676
rect 27105 4642 27114 4676
rect 27062 4633 27114 4642
rect 26972 4388 27024 4391
rect 26972 4354 26981 4388
rect 26981 4354 27015 4388
rect 27015 4354 27024 4388
rect 26972 4339 27024 4354
rect 27152 4388 27204 4391
rect 27152 4354 27161 4388
rect 27161 4354 27195 4388
rect 27195 4354 27204 4388
rect 27152 4339 27204 4354
rect 15380 4243 15432 4295
rect 15560 4243 15612 4295
rect 15819 4243 15871 4295
rect 15883 4243 15935 4295
rect 26972 4243 27024 4295
rect 27152 4243 27204 4295
rect 27411 4243 27463 4295
rect 27475 4243 27527 4295
rect 12897 4065 12949 4117
rect 13396 4065 13448 4117
rect 13786 4065 13838 4117
rect 14176 4065 14228 4117
rect 14566 4065 14618 4117
rect 14956 4065 15008 4117
rect 15671 4065 15723 4117
rect 24489 4065 24541 4117
rect 24988 4065 25040 4117
rect 25378 4065 25430 4117
rect 25768 4065 25820 4117
rect 26158 4065 26210 4117
rect 26548 4065 26600 4117
rect 27263 4065 27315 4117
rect 12596 3908 12648 3960
rect 24188 3908 24240 3960
rect 13006 3472 13058 3477
rect 13006 3438 13015 3472
rect 13015 3438 13049 3472
rect 13049 3438 13058 3472
rect 13006 3425 13058 3438
rect 12596 3346 12648 3398
rect 13006 3400 13058 3413
rect 13006 3366 13015 3400
rect 13015 3366 13049 3400
rect 13049 3366 13058 3400
rect 13006 3361 13058 3366
rect 13396 3820 13448 3825
rect 13396 3786 13405 3820
rect 13405 3786 13439 3820
rect 13439 3786 13448 3820
rect 13396 3773 13448 3786
rect 13396 3748 13448 3761
rect 13396 3714 13405 3748
rect 13405 3714 13439 3748
rect 13439 3714 13448 3748
rect 13396 3709 13448 3714
rect 13526 3820 13578 3825
rect 13526 3786 13535 3820
rect 13535 3786 13569 3820
rect 13569 3786 13578 3820
rect 13526 3773 13578 3786
rect 13526 3748 13578 3761
rect 13526 3714 13535 3748
rect 13535 3714 13569 3748
rect 13569 3714 13578 3748
rect 13526 3709 13578 3714
rect 13136 3438 13145 3445
rect 13145 3438 13179 3445
rect 13179 3438 13188 3445
rect 13136 3400 13188 3438
rect 13136 3393 13145 3400
rect 13145 3393 13179 3400
rect 13179 3393 13188 3400
rect 13396 3438 13405 3445
rect 13405 3438 13439 3445
rect 13439 3438 13448 3445
rect 13396 3400 13448 3438
rect 13396 3393 13405 3400
rect 13405 3393 13439 3400
rect 13439 3393 13448 3400
rect 13786 3820 13838 3825
rect 13786 3786 13795 3820
rect 13795 3786 13829 3820
rect 13829 3786 13838 3820
rect 13786 3773 13838 3786
rect 13786 3748 13838 3761
rect 13786 3714 13795 3748
rect 13795 3714 13829 3748
rect 13829 3714 13838 3748
rect 13786 3709 13838 3714
rect 13916 3820 13968 3825
rect 13916 3786 13925 3820
rect 13925 3786 13959 3820
rect 13959 3786 13968 3820
rect 13916 3773 13968 3786
rect 13916 3748 13968 3761
rect 13916 3714 13925 3748
rect 13925 3714 13959 3748
rect 13959 3714 13968 3748
rect 13916 3709 13968 3714
rect 13526 3438 13535 3445
rect 13535 3438 13569 3445
rect 13569 3438 13578 3445
rect 13526 3400 13578 3438
rect 13526 3393 13535 3400
rect 13535 3393 13569 3400
rect 13569 3393 13578 3400
rect 13786 3438 13795 3445
rect 13795 3438 13829 3445
rect 13829 3438 13838 3445
rect 13786 3400 13838 3438
rect 13786 3393 13795 3400
rect 13795 3393 13829 3400
rect 13829 3393 13838 3400
rect 14176 3820 14228 3825
rect 14176 3786 14185 3820
rect 14185 3786 14219 3820
rect 14219 3786 14228 3820
rect 14176 3773 14228 3786
rect 14176 3748 14228 3761
rect 14176 3714 14185 3748
rect 14185 3714 14219 3748
rect 14219 3714 14228 3748
rect 14176 3709 14228 3714
rect 14306 3820 14358 3825
rect 14306 3786 14315 3820
rect 14315 3786 14349 3820
rect 14349 3786 14358 3820
rect 14306 3773 14358 3786
rect 14306 3748 14358 3761
rect 14306 3714 14315 3748
rect 14315 3714 14349 3748
rect 14349 3714 14358 3748
rect 14306 3709 14358 3714
rect 13916 3438 13925 3445
rect 13925 3438 13959 3445
rect 13959 3438 13968 3445
rect 13916 3400 13968 3438
rect 13916 3393 13925 3400
rect 13925 3393 13959 3400
rect 13959 3393 13968 3400
rect 14176 3438 14185 3445
rect 14185 3438 14219 3445
rect 14219 3438 14228 3445
rect 14176 3400 14228 3438
rect 14176 3393 14185 3400
rect 14185 3393 14219 3400
rect 14219 3393 14228 3400
rect 14566 3820 14618 3825
rect 14566 3786 14575 3820
rect 14575 3786 14609 3820
rect 14609 3786 14618 3820
rect 14566 3773 14618 3786
rect 14566 3748 14618 3761
rect 14566 3714 14575 3748
rect 14575 3714 14609 3748
rect 14609 3714 14618 3748
rect 14566 3709 14618 3714
rect 14696 3820 14748 3825
rect 14696 3786 14705 3820
rect 14705 3786 14739 3820
rect 14739 3786 14748 3820
rect 14696 3773 14748 3786
rect 14696 3748 14748 3761
rect 14696 3714 14705 3748
rect 14705 3714 14739 3748
rect 14739 3714 14748 3748
rect 14696 3709 14748 3714
rect 14306 3438 14315 3445
rect 14315 3438 14349 3445
rect 14349 3438 14358 3445
rect 14306 3400 14358 3438
rect 14306 3393 14315 3400
rect 14315 3393 14349 3400
rect 14349 3393 14358 3400
rect 14566 3438 14575 3445
rect 14575 3438 14609 3445
rect 14609 3438 14618 3445
rect 14566 3400 14618 3438
rect 14566 3393 14575 3400
rect 14575 3393 14609 3400
rect 14609 3393 14618 3400
rect 14956 3820 15008 3825
rect 14956 3786 14965 3820
rect 14965 3786 14999 3820
rect 14999 3786 15008 3820
rect 14956 3773 15008 3786
rect 14956 3748 15008 3761
rect 14956 3714 14965 3748
rect 14965 3714 14999 3748
rect 14999 3714 15008 3748
rect 14956 3709 15008 3714
rect 15086 3820 15138 3825
rect 15086 3786 15095 3820
rect 15095 3786 15129 3820
rect 15129 3786 15138 3820
rect 15086 3773 15138 3786
rect 15200 3820 15252 3829
rect 15200 3786 15209 3820
rect 15209 3786 15243 3820
rect 15243 3786 15252 3820
rect 15200 3777 15252 3786
rect 15086 3748 15138 3761
rect 15086 3714 15095 3748
rect 15095 3714 15129 3748
rect 15129 3714 15138 3748
rect 15086 3709 15138 3714
rect 15380 3820 15432 3829
rect 15380 3786 15389 3820
rect 15389 3786 15423 3820
rect 15423 3786 15432 3820
rect 15380 3777 15432 3786
rect 15290 3748 15342 3757
rect 15290 3714 15299 3748
rect 15299 3714 15333 3748
rect 15333 3714 15342 3748
rect 15290 3705 15342 3714
rect 15560 3820 15612 3829
rect 15560 3786 15569 3820
rect 15569 3786 15603 3820
rect 15603 3786 15612 3820
rect 15560 3777 15612 3786
rect 15470 3748 15522 3757
rect 15470 3714 15479 3748
rect 15479 3714 15513 3748
rect 15513 3714 15522 3748
rect 15470 3705 15522 3714
rect 15316 3579 15368 3588
rect 15316 3545 15318 3579
rect 15318 3545 15352 3579
rect 15352 3545 15368 3579
rect 15316 3536 15368 3545
rect 15380 3579 15432 3588
rect 15380 3545 15390 3579
rect 15390 3545 15424 3579
rect 15424 3545 15432 3579
rect 15380 3536 15432 3545
rect 15444 3579 15496 3588
rect 15444 3545 15462 3579
rect 15462 3545 15496 3579
rect 15444 3536 15496 3545
rect 14696 3438 14705 3445
rect 14705 3438 14739 3445
rect 14739 3438 14748 3445
rect 14696 3400 14748 3438
rect 14696 3393 14705 3400
rect 14705 3393 14739 3400
rect 14739 3393 14748 3400
rect 14956 3438 14965 3445
rect 14965 3438 14999 3445
rect 14999 3438 15008 3445
rect 14956 3400 15008 3438
rect 14956 3393 14965 3400
rect 14965 3393 14999 3400
rect 14999 3393 15008 3400
rect 15086 3438 15095 3445
rect 15095 3438 15129 3445
rect 15129 3438 15138 3445
rect 15086 3400 15138 3438
rect 15086 3393 15095 3400
rect 15095 3393 15129 3400
rect 15129 3393 15138 3400
rect 24598 3472 24650 3477
rect 24598 3438 24607 3472
rect 24607 3438 24641 3472
rect 24641 3438 24650 3472
rect 24598 3425 24650 3438
rect 24188 3346 24240 3398
rect 24598 3400 24650 3413
rect 24598 3366 24607 3400
rect 24607 3366 24641 3400
rect 24641 3366 24650 3400
rect 24598 3361 24650 3366
rect 24988 3820 25040 3825
rect 24988 3786 24997 3820
rect 24997 3786 25031 3820
rect 25031 3786 25040 3820
rect 24988 3773 25040 3786
rect 24988 3748 25040 3761
rect 24988 3714 24997 3748
rect 24997 3714 25031 3748
rect 25031 3714 25040 3748
rect 24988 3709 25040 3714
rect 25118 3820 25170 3825
rect 25118 3786 25127 3820
rect 25127 3786 25161 3820
rect 25161 3786 25170 3820
rect 25118 3773 25170 3786
rect 25118 3748 25170 3761
rect 25118 3714 25127 3748
rect 25127 3714 25161 3748
rect 25161 3714 25170 3748
rect 25118 3709 25170 3714
rect 24728 3438 24737 3445
rect 24737 3438 24771 3445
rect 24771 3438 24780 3445
rect 24728 3400 24780 3438
rect 24728 3393 24737 3400
rect 24737 3393 24771 3400
rect 24771 3393 24780 3400
rect 24988 3438 24997 3445
rect 24997 3438 25031 3445
rect 25031 3438 25040 3445
rect 24988 3400 25040 3438
rect 24988 3393 24997 3400
rect 24997 3393 25031 3400
rect 25031 3393 25040 3400
rect 25378 3820 25430 3825
rect 25378 3786 25387 3820
rect 25387 3786 25421 3820
rect 25421 3786 25430 3820
rect 25378 3773 25430 3786
rect 25378 3748 25430 3761
rect 25378 3714 25387 3748
rect 25387 3714 25421 3748
rect 25421 3714 25430 3748
rect 25378 3709 25430 3714
rect 25508 3820 25560 3825
rect 25508 3786 25517 3820
rect 25517 3786 25551 3820
rect 25551 3786 25560 3820
rect 25508 3773 25560 3786
rect 25508 3748 25560 3761
rect 25508 3714 25517 3748
rect 25517 3714 25551 3748
rect 25551 3714 25560 3748
rect 25508 3709 25560 3714
rect 25118 3438 25127 3445
rect 25127 3438 25161 3445
rect 25161 3438 25170 3445
rect 25118 3400 25170 3438
rect 25118 3393 25127 3400
rect 25127 3393 25161 3400
rect 25161 3393 25170 3400
rect 25378 3438 25387 3445
rect 25387 3438 25421 3445
rect 25421 3438 25430 3445
rect 25378 3400 25430 3438
rect 25378 3393 25387 3400
rect 25387 3393 25421 3400
rect 25421 3393 25430 3400
rect 25768 3820 25820 3825
rect 25768 3786 25777 3820
rect 25777 3786 25811 3820
rect 25811 3786 25820 3820
rect 25768 3773 25820 3786
rect 25768 3748 25820 3761
rect 25768 3714 25777 3748
rect 25777 3714 25811 3748
rect 25811 3714 25820 3748
rect 25768 3709 25820 3714
rect 25898 3820 25950 3825
rect 25898 3786 25907 3820
rect 25907 3786 25941 3820
rect 25941 3786 25950 3820
rect 25898 3773 25950 3786
rect 25898 3748 25950 3761
rect 25898 3714 25907 3748
rect 25907 3714 25941 3748
rect 25941 3714 25950 3748
rect 25898 3709 25950 3714
rect 25508 3438 25517 3445
rect 25517 3438 25551 3445
rect 25551 3438 25560 3445
rect 25508 3400 25560 3438
rect 25508 3393 25517 3400
rect 25517 3393 25551 3400
rect 25551 3393 25560 3400
rect 25768 3438 25777 3445
rect 25777 3438 25811 3445
rect 25811 3438 25820 3445
rect 25768 3400 25820 3438
rect 25768 3393 25777 3400
rect 25777 3393 25811 3400
rect 25811 3393 25820 3400
rect 26158 3820 26210 3825
rect 26158 3786 26167 3820
rect 26167 3786 26201 3820
rect 26201 3786 26210 3820
rect 26158 3773 26210 3786
rect 26158 3748 26210 3761
rect 26158 3714 26167 3748
rect 26167 3714 26201 3748
rect 26201 3714 26210 3748
rect 26158 3709 26210 3714
rect 26288 3820 26340 3825
rect 26288 3786 26297 3820
rect 26297 3786 26331 3820
rect 26331 3786 26340 3820
rect 26288 3773 26340 3786
rect 26288 3748 26340 3761
rect 26288 3714 26297 3748
rect 26297 3714 26331 3748
rect 26331 3714 26340 3748
rect 26288 3709 26340 3714
rect 25898 3438 25907 3445
rect 25907 3438 25941 3445
rect 25941 3438 25950 3445
rect 25898 3400 25950 3438
rect 25898 3393 25907 3400
rect 25907 3393 25941 3400
rect 25941 3393 25950 3400
rect 26158 3438 26167 3445
rect 26167 3438 26201 3445
rect 26201 3438 26210 3445
rect 26158 3400 26210 3438
rect 26158 3393 26167 3400
rect 26167 3393 26201 3400
rect 26201 3393 26210 3400
rect 26548 3820 26600 3825
rect 26548 3786 26557 3820
rect 26557 3786 26591 3820
rect 26591 3786 26600 3820
rect 26548 3773 26600 3786
rect 26548 3748 26600 3761
rect 26548 3714 26557 3748
rect 26557 3714 26591 3748
rect 26591 3714 26600 3748
rect 26548 3709 26600 3714
rect 26678 3820 26730 3825
rect 26678 3786 26687 3820
rect 26687 3786 26721 3820
rect 26721 3786 26730 3820
rect 26678 3773 26730 3786
rect 26792 3820 26844 3829
rect 26792 3786 26801 3820
rect 26801 3786 26835 3820
rect 26835 3786 26844 3820
rect 26792 3777 26844 3786
rect 26678 3748 26730 3761
rect 26678 3714 26687 3748
rect 26687 3714 26721 3748
rect 26721 3714 26730 3748
rect 26678 3709 26730 3714
rect 26972 3820 27024 3829
rect 26972 3786 26981 3820
rect 26981 3786 27015 3820
rect 27015 3786 27024 3820
rect 26972 3777 27024 3786
rect 26882 3748 26934 3757
rect 26882 3714 26891 3748
rect 26891 3714 26925 3748
rect 26925 3714 26934 3748
rect 26882 3705 26934 3714
rect 27152 3820 27204 3829
rect 27152 3786 27161 3820
rect 27161 3786 27195 3820
rect 27195 3786 27204 3820
rect 27152 3777 27204 3786
rect 27062 3748 27114 3757
rect 27062 3714 27071 3748
rect 27071 3714 27105 3748
rect 27105 3714 27114 3748
rect 27062 3705 27114 3714
rect 26908 3579 26960 3588
rect 26908 3545 26910 3579
rect 26910 3545 26944 3579
rect 26944 3545 26960 3579
rect 26908 3536 26960 3545
rect 26972 3579 27024 3588
rect 26972 3545 26982 3579
rect 26982 3545 27016 3579
rect 27016 3545 27024 3579
rect 26972 3536 27024 3545
rect 27036 3579 27088 3588
rect 27036 3545 27054 3579
rect 27054 3545 27088 3579
rect 27036 3536 27088 3545
rect 26288 3438 26297 3445
rect 26297 3438 26331 3445
rect 26331 3438 26340 3445
rect 26288 3400 26340 3438
rect 26288 3393 26297 3400
rect 26297 3393 26331 3400
rect 26331 3393 26340 3400
rect 26548 3438 26557 3445
rect 26557 3438 26591 3445
rect 26591 3438 26600 3445
rect 26548 3400 26600 3438
rect 26548 3393 26557 3400
rect 26557 3393 26591 3400
rect 26591 3393 26600 3400
rect 26678 3438 26687 3445
rect 26687 3438 26721 3445
rect 26721 3438 26730 3445
rect 26678 3400 26730 3438
rect 26678 3393 26687 3400
rect 26687 3393 26721 3400
rect 26721 3393 26730 3400
rect 12688 3220 12740 3272
rect 13003 3263 13055 3272
rect 13003 3229 13012 3263
rect 13012 3229 13046 3263
rect 13046 3229 13055 3263
rect 13003 3220 13055 3229
rect 13331 3263 13383 3272
rect 13331 3229 13340 3263
rect 13340 3229 13374 3263
rect 13374 3229 13383 3263
rect 13331 3220 13383 3229
rect 13721 3263 13773 3272
rect 13721 3229 13730 3263
rect 13730 3229 13764 3263
rect 13764 3229 13773 3263
rect 13721 3220 13773 3229
rect 14111 3263 14163 3272
rect 14111 3229 14120 3263
rect 14120 3229 14154 3263
rect 14154 3229 14163 3263
rect 14111 3220 14163 3229
rect 14501 3263 14553 3272
rect 14501 3229 14510 3263
rect 14510 3229 14544 3263
rect 14544 3229 14553 3263
rect 14501 3220 14553 3229
rect 14891 3263 14943 3272
rect 14891 3229 14900 3263
rect 14900 3229 14934 3263
rect 14934 3229 14943 3263
rect 14891 3220 14943 3229
rect 24280 3220 24332 3272
rect 24595 3263 24647 3272
rect 24595 3229 24604 3263
rect 24604 3229 24638 3263
rect 24638 3229 24647 3263
rect 24595 3220 24647 3229
rect 24923 3263 24975 3272
rect 24923 3229 24932 3263
rect 24932 3229 24966 3263
rect 24966 3229 24975 3263
rect 24923 3220 24975 3229
rect 25313 3263 25365 3272
rect 25313 3229 25322 3263
rect 25322 3229 25356 3263
rect 25356 3229 25365 3263
rect 25313 3220 25365 3229
rect 25703 3263 25755 3272
rect 25703 3229 25712 3263
rect 25712 3229 25746 3263
rect 25746 3229 25755 3263
rect 25703 3220 25755 3229
rect 26093 3263 26145 3272
rect 26093 3229 26102 3263
rect 26102 3229 26136 3263
rect 26136 3229 26145 3263
rect 26093 3220 26145 3229
rect 26483 3263 26535 3272
rect 26483 3229 26492 3263
rect 26492 3229 26526 3263
rect 26526 3229 26535 3263
rect 26483 3220 26535 3229
rect 13267 3130 13319 3139
rect 13267 3096 13268 3130
rect 13268 3096 13302 3130
rect 13302 3096 13319 3130
rect 13267 3087 13319 3096
rect 13331 3130 13383 3139
rect 13331 3096 13340 3130
rect 13340 3096 13374 3130
rect 13374 3096 13383 3130
rect 13331 3087 13383 3096
rect 13395 3130 13447 3139
rect 14047 3130 14099 3139
rect 13395 3096 13412 3130
rect 13412 3096 13446 3130
rect 13446 3096 13447 3130
rect 14047 3096 14048 3130
rect 14048 3096 14082 3130
rect 14082 3096 14099 3130
rect 13395 3087 13447 3096
rect 14047 3087 14099 3096
rect 14111 3130 14163 3139
rect 14111 3096 14120 3130
rect 14120 3096 14154 3130
rect 14154 3096 14163 3130
rect 14111 3087 14163 3096
rect 14175 3130 14227 3139
rect 14827 3130 14879 3139
rect 14175 3096 14192 3130
rect 14192 3096 14226 3130
rect 14226 3096 14227 3130
rect 14827 3096 14828 3130
rect 14828 3096 14862 3130
rect 14862 3096 14879 3130
rect 14175 3087 14227 3096
rect 14827 3087 14879 3096
rect 14891 3130 14943 3139
rect 14891 3096 14900 3130
rect 14900 3096 14934 3130
rect 14934 3096 14943 3130
rect 14891 3087 14943 3096
rect 14955 3130 15007 3139
rect 14955 3096 14972 3130
rect 14972 3096 15006 3130
rect 15006 3096 15007 3130
rect 14955 3087 15007 3096
rect 24859 3130 24911 3139
rect 24859 3096 24860 3130
rect 24860 3096 24894 3130
rect 24894 3096 24911 3130
rect 24859 3087 24911 3096
rect 24923 3130 24975 3139
rect 24923 3096 24932 3130
rect 24932 3096 24966 3130
rect 24966 3096 24975 3130
rect 24923 3087 24975 3096
rect 24987 3130 25039 3139
rect 25639 3130 25691 3139
rect 24987 3096 25004 3130
rect 25004 3096 25038 3130
rect 25038 3096 25039 3130
rect 25639 3096 25640 3130
rect 25640 3096 25674 3130
rect 25674 3096 25691 3130
rect 24987 3087 25039 3096
rect 25639 3087 25691 3096
rect 25703 3130 25755 3139
rect 25703 3096 25712 3130
rect 25712 3096 25746 3130
rect 25746 3096 25755 3130
rect 25703 3087 25755 3096
rect 25767 3130 25819 3139
rect 26419 3130 26471 3139
rect 25767 3096 25784 3130
rect 25784 3096 25818 3130
rect 25818 3096 25819 3130
rect 26419 3096 26420 3130
rect 26420 3096 26454 3130
rect 26454 3096 26471 3130
rect 25767 3087 25819 3096
rect 26419 3087 26471 3096
rect 26483 3130 26535 3139
rect 26483 3096 26492 3130
rect 26492 3096 26526 3130
rect 26526 3096 26535 3130
rect 26483 3087 26535 3096
rect 26547 3130 26599 3139
rect 26547 3096 26564 3130
rect 26564 3096 26598 3130
rect 26598 3096 26599 3130
rect 26547 3087 26599 3096
rect 12688 2954 12740 3006
rect 13331 2997 13383 3006
rect 13331 2963 13340 2997
rect 13340 2963 13374 2997
rect 13374 2963 13383 2997
rect 13331 2954 13383 2963
rect 13721 2997 13773 3006
rect 13721 2963 13730 2997
rect 13730 2963 13764 2997
rect 13764 2963 13773 2997
rect 13721 2954 13773 2963
rect 14111 2997 14163 3006
rect 14111 2963 14120 2997
rect 14120 2963 14154 2997
rect 14154 2963 14163 2997
rect 14111 2954 14163 2963
rect 14501 2997 14553 3006
rect 14501 2963 14510 2997
rect 14510 2963 14544 2997
rect 14544 2963 14553 2997
rect 14501 2954 14553 2963
rect 14891 2997 14943 3006
rect 14891 2963 14900 2997
rect 14900 2963 14934 2997
rect 14934 2963 14943 2997
rect 14891 2954 14943 2963
rect 15281 2997 15333 3006
rect 15281 2963 15290 2997
rect 15290 2963 15324 2997
rect 15324 2963 15333 2997
rect 15281 2954 15333 2963
rect 24280 2954 24332 3006
rect 24923 2997 24975 3006
rect 24923 2963 24932 2997
rect 24932 2963 24966 2997
rect 24966 2963 24975 2997
rect 24923 2954 24975 2963
rect 25313 2997 25365 3006
rect 25313 2963 25322 2997
rect 25322 2963 25356 2997
rect 25356 2963 25365 2997
rect 25313 2954 25365 2963
rect 25703 2997 25755 3006
rect 25703 2963 25712 2997
rect 25712 2963 25746 2997
rect 25746 2963 25755 2997
rect 25703 2954 25755 2963
rect 26093 2997 26145 3006
rect 26093 2963 26102 2997
rect 26102 2963 26136 2997
rect 26136 2963 26145 2997
rect 26093 2954 26145 2963
rect 26483 2997 26535 3006
rect 26483 2963 26492 2997
rect 26492 2963 26526 2997
rect 26526 2963 26535 2997
rect 26483 2954 26535 2963
rect 26873 2997 26925 3006
rect 26873 2963 26882 2997
rect 26882 2963 26916 2997
rect 26916 2963 26925 2997
rect 26873 2954 26925 2963
rect 13136 2826 13145 2833
rect 13145 2826 13179 2833
rect 13179 2826 13188 2833
rect 13136 2788 13188 2826
rect 13136 2781 13145 2788
rect 13145 2781 13179 2788
rect 13179 2781 13188 2788
rect 13266 2826 13275 2833
rect 13275 2826 13309 2833
rect 13309 2826 13318 2833
rect 13266 2788 13318 2826
rect 13266 2781 13275 2788
rect 13275 2781 13309 2788
rect 13309 2781 13318 2788
rect 13526 2826 13535 2833
rect 13535 2826 13569 2833
rect 13569 2826 13578 2833
rect 13526 2788 13578 2826
rect 13526 2781 13535 2788
rect 13535 2781 13569 2788
rect 13569 2781 13578 2788
rect 13136 2512 13188 2517
rect 13136 2478 13145 2512
rect 13145 2478 13179 2512
rect 13179 2478 13188 2512
rect 13136 2465 13188 2478
rect 13136 2440 13188 2453
rect 13136 2406 13145 2440
rect 13145 2406 13179 2440
rect 13179 2406 13188 2440
rect 13136 2401 13188 2406
rect 13266 2512 13318 2517
rect 13266 2478 13275 2512
rect 13275 2478 13309 2512
rect 13309 2478 13318 2512
rect 13266 2465 13318 2478
rect 13266 2440 13318 2453
rect 13266 2406 13275 2440
rect 13275 2406 13309 2440
rect 13309 2406 13318 2440
rect 13266 2401 13318 2406
rect 13656 2826 13665 2833
rect 13665 2826 13699 2833
rect 13699 2826 13708 2833
rect 13656 2788 13708 2826
rect 13656 2781 13665 2788
rect 13665 2781 13699 2788
rect 13699 2781 13708 2788
rect 13916 2826 13925 2833
rect 13925 2826 13959 2833
rect 13959 2826 13968 2833
rect 13916 2788 13968 2826
rect 13916 2781 13925 2788
rect 13925 2781 13959 2788
rect 13959 2781 13968 2788
rect 13526 2512 13578 2517
rect 13526 2478 13535 2512
rect 13535 2478 13569 2512
rect 13569 2478 13578 2512
rect 13526 2465 13578 2478
rect 13526 2440 13578 2453
rect 13526 2406 13535 2440
rect 13535 2406 13569 2440
rect 13569 2406 13578 2440
rect 13526 2401 13578 2406
rect 13656 2512 13708 2517
rect 13656 2478 13665 2512
rect 13665 2478 13699 2512
rect 13699 2478 13708 2512
rect 13656 2465 13708 2478
rect 13656 2440 13708 2453
rect 13656 2406 13665 2440
rect 13665 2406 13699 2440
rect 13699 2406 13708 2440
rect 13656 2401 13708 2406
rect 14046 2826 14055 2833
rect 14055 2826 14089 2833
rect 14089 2826 14098 2833
rect 14046 2788 14098 2826
rect 14046 2781 14055 2788
rect 14055 2781 14089 2788
rect 14089 2781 14098 2788
rect 14306 2826 14315 2833
rect 14315 2826 14349 2833
rect 14349 2826 14358 2833
rect 14306 2788 14358 2826
rect 14306 2781 14315 2788
rect 14315 2781 14349 2788
rect 14349 2781 14358 2788
rect 13916 2512 13968 2517
rect 13916 2478 13925 2512
rect 13925 2478 13959 2512
rect 13959 2478 13968 2512
rect 13916 2465 13968 2478
rect 13916 2440 13968 2453
rect 13916 2406 13925 2440
rect 13925 2406 13959 2440
rect 13959 2406 13968 2440
rect 13916 2401 13968 2406
rect 14046 2512 14098 2517
rect 14046 2478 14055 2512
rect 14055 2478 14089 2512
rect 14089 2478 14098 2512
rect 14046 2465 14098 2478
rect 14046 2440 14098 2453
rect 14046 2406 14055 2440
rect 14055 2406 14089 2440
rect 14089 2406 14098 2440
rect 14046 2401 14098 2406
rect 14436 2826 14445 2833
rect 14445 2826 14479 2833
rect 14479 2826 14488 2833
rect 14436 2788 14488 2826
rect 14436 2781 14445 2788
rect 14445 2781 14479 2788
rect 14479 2781 14488 2788
rect 14696 2826 14705 2833
rect 14705 2826 14739 2833
rect 14739 2826 14748 2833
rect 14696 2788 14748 2826
rect 14696 2781 14705 2788
rect 14705 2781 14739 2788
rect 14739 2781 14748 2788
rect 14306 2512 14358 2517
rect 14306 2478 14315 2512
rect 14315 2478 14349 2512
rect 14349 2478 14358 2512
rect 14306 2465 14358 2478
rect 14306 2440 14358 2453
rect 14306 2406 14315 2440
rect 14315 2406 14349 2440
rect 14349 2406 14358 2440
rect 14306 2401 14358 2406
rect 14436 2512 14488 2517
rect 14436 2478 14445 2512
rect 14445 2478 14479 2512
rect 14479 2478 14488 2512
rect 14436 2465 14488 2478
rect 14436 2440 14488 2453
rect 14436 2406 14445 2440
rect 14445 2406 14479 2440
rect 14479 2406 14488 2440
rect 14436 2401 14488 2406
rect 14826 2826 14835 2833
rect 14835 2826 14869 2833
rect 14869 2826 14878 2833
rect 14826 2788 14878 2826
rect 14826 2781 14835 2788
rect 14835 2781 14869 2788
rect 14869 2781 14878 2788
rect 15086 2826 15095 2833
rect 15095 2826 15129 2833
rect 15129 2826 15138 2833
rect 15086 2788 15138 2826
rect 15086 2781 15095 2788
rect 15095 2781 15129 2788
rect 15129 2781 15138 2788
rect 14696 2512 14748 2517
rect 14696 2478 14705 2512
rect 14705 2478 14739 2512
rect 14739 2478 14748 2512
rect 14696 2465 14748 2478
rect 14696 2440 14748 2453
rect 14696 2406 14705 2440
rect 14705 2406 14739 2440
rect 14739 2406 14748 2440
rect 14696 2401 14748 2406
rect 14826 2512 14878 2517
rect 14826 2478 14835 2512
rect 14835 2478 14869 2512
rect 14869 2478 14878 2512
rect 14826 2465 14878 2478
rect 14826 2440 14878 2453
rect 14826 2406 14835 2440
rect 14835 2406 14869 2440
rect 14869 2406 14878 2440
rect 14826 2401 14878 2406
rect 15216 2826 15225 2833
rect 15225 2826 15259 2833
rect 15259 2826 15268 2833
rect 15216 2788 15268 2826
rect 15216 2781 15225 2788
rect 15225 2781 15259 2788
rect 15259 2781 15268 2788
rect 15476 2826 15485 2833
rect 15485 2826 15519 2833
rect 15519 2826 15528 2833
rect 15476 2788 15528 2826
rect 15476 2781 15485 2788
rect 15485 2781 15519 2788
rect 15519 2781 15528 2788
rect 15086 2512 15138 2517
rect 15086 2478 15095 2512
rect 15095 2478 15129 2512
rect 15129 2478 15138 2512
rect 15086 2465 15138 2478
rect 15086 2440 15138 2453
rect 15086 2406 15095 2440
rect 15095 2406 15129 2440
rect 15129 2406 15138 2440
rect 15086 2401 15138 2406
rect 15216 2512 15268 2517
rect 15216 2478 15225 2512
rect 15225 2478 15259 2512
rect 15259 2478 15268 2512
rect 15216 2465 15268 2478
rect 15216 2440 15268 2453
rect 15216 2406 15225 2440
rect 15225 2406 15259 2440
rect 15259 2406 15268 2440
rect 15216 2401 15268 2406
rect 24728 2826 24737 2833
rect 24737 2826 24771 2833
rect 24771 2826 24780 2833
rect 24728 2788 24780 2826
rect 24728 2781 24737 2788
rect 24737 2781 24771 2788
rect 24771 2781 24780 2788
rect 24858 2826 24867 2833
rect 24867 2826 24901 2833
rect 24901 2826 24910 2833
rect 24858 2788 24910 2826
rect 24858 2781 24867 2788
rect 24867 2781 24901 2788
rect 24901 2781 24910 2788
rect 25118 2826 25127 2833
rect 25127 2826 25161 2833
rect 25161 2826 25170 2833
rect 25118 2788 25170 2826
rect 25118 2781 25127 2788
rect 25127 2781 25161 2788
rect 25161 2781 25170 2788
rect 24728 2512 24780 2517
rect 24728 2478 24737 2512
rect 24737 2478 24771 2512
rect 24771 2478 24780 2512
rect 24728 2465 24780 2478
rect 24728 2440 24780 2453
rect 24728 2406 24737 2440
rect 24737 2406 24771 2440
rect 24771 2406 24780 2440
rect 24728 2401 24780 2406
rect 24858 2512 24910 2517
rect 24858 2478 24867 2512
rect 24867 2478 24901 2512
rect 24901 2478 24910 2512
rect 24858 2465 24910 2478
rect 24858 2440 24910 2453
rect 24858 2406 24867 2440
rect 24867 2406 24901 2440
rect 24901 2406 24910 2440
rect 24858 2401 24910 2406
rect 25248 2826 25257 2833
rect 25257 2826 25291 2833
rect 25291 2826 25300 2833
rect 25248 2788 25300 2826
rect 25248 2781 25257 2788
rect 25257 2781 25291 2788
rect 25291 2781 25300 2788
rect 25508 2826 25517 2833
rect 25517 2826 25551 2833
rect 25551 2826 25560 2833
rect 25508 2788 25560 2826
rect 25508 2781 25517 2788
rect 25517 2781 25551 2788
rect 25551 2781 25560 2788
rect 25118 2512 25170 2517
rect 25118 2478 25127 2512
rect 25127 2478 25161 2512
rect 25161 2478 25170 2512
rect 25118 2465 25170 2478
rect 25118 2440 25170 2453
rect 25118 2406 25127 2440
rect 25127 2406 25161 2440
rect 25161 2406 25170 2440
rect 25118 2401 25170 2406
rect 25248 2512 25300 2517
rect 25248 2478 25257 2512
rect 25257 2478 25291 2512
rect 25291 2478 25300 2512
rect 25248 2465 25300 2478
rect 25248 2440 25300 2453
rect 25248 2406 25257 2440
rect 25257 2406 25291 2440
rect 25291 2406 25300 2440
rect 25248 2401 25300 2406
rect 25638 2826 25647 2833
rect 25647 2826 25681 2833
rect 25681 2826 25690 2833
rect 25638 2788 25690 2826
rect 25638 2781 25647 2788
rect 25647 2781 25681 2788
rect 25681 2781 25690 2788
rect 25898 2826 25907 2833
rect 25907 2826 25941 2833
rect 25941 2826 25950 2833
rect 25898 2788 25950 2826
rect 25898 2781 25907 2788
rect 25907 2781 25941 2788
rect 25941 2781 25950 2788
rect 25508 2512 25560 2517
rect 25508 2478 25517 2512
rect 25517 2478 25551 2512
rect 25551 2478 25560 2512
rect 25508 2465 25560 2478
rect 25508 2440 25560 2453
rect 25508 2406 25517 2440
rect 25517 2406 25551 2440
rect 25551 2406 25560 2440
rect 25508 2401 25560 2406
rect 25638 2512 25690 2517
rect 25638 2478 25647 2512
rect 25647 2478 25681 2512
rect 25681 2478 25690 2512
rect 25638 2465 25690 2478
rect 25638 2440 25690 2453
rect 25638 2406 25647 2440
rect 25647 2406 25681 2440
rect 25681 2406 25690 2440
rect 25638 2401 25690 2406
rect 26028 2826 26037 2833
rect 26037 2826 26071 2833
rect 26071 2826 26080 2833
rect 26028 2788 26080 2826
rect 26028 2781 26037 2788
rect 26037 2781 26071 2788
rect 26071 2781 26080 2788
rect 26288 2826 26297 2833
rect 26297 2826 26331 2833
rect 26331 2826 26340 2833
rect 26288 2788 26340 2826
rect 26288 2781 26297 2788
rect 26297 2781 26331 2788
rect 26331 2781 26340 2788
rect 25898 2512 25950 2517
rect 25898 2478 25907 2512
rect 25907 2478 25941 2512
rect 25941 2478 25950 2512
rect 25898 2465 25950 2478
rect 25898 2440 25950 2453
rect 25898 2406 25907 2440
rect 25907 2406 25941 2440
rect 25941 2406 25950 2440
rect 25898 2401 25950 2406
rect 26028 2512 26080 2517
rect 26028 2478 26037 2512
rect 26037 2478 26071 2512
rect 26071 2478 26080 2512
rect 26028 2465 26080 2478
rect 26028 2440 26080 2453
rect 26028 2406 26037 2440
rect 26037 2406 26071 2440
rect 26071 2406 26080 2440
rect 26028 2401 26080 2406
rect 26418 2826 26427 2833
rect 26427 2826 26461 2833
rect 26461 2826 26470 2833
rect 26418 2788 26470 2826
rect 26418 2781 26427 2788
rect 26427 2781 26461 2788
rect 26461 2781 26470 2788
rect 26678 2826 26687 2833
rect 26687 2826 26721 2833
rect 26721 2826 26730 2833
rect 26678 2788 26730 2826
rect 26678 2781 26687 2788
rect 26687 2781 26721 2788
rect 26721 2781 26730 2788
rect 26288 2512 26340 2517
rect 26288 2478 26297 2512
rect 26297 2478 26331 2512
rect 26331 2478 26340 2512
rect 26288 2465 26340 2478
rect 26288 2440 26340 2453
rect 26288 2406 26297 2440
rect 26297 2406 26331 2440
rect 26331 2406 26340 2440
rect 26288 2401 26340 2406
rect 26418 2512 26470 2517
rect 26418 2478 26427 2512
rect 26427 2478 26461 2512
rect 26461 2478 26470 2512
rect 26418 2465 26470 2478
rect 26418 2440 26470 2453
rect 26418 2406 26427 2440
rect 26427 2406 26461 2440
rect 26461 2406 26470 2440
rect 26418 2401 26470 2406
rect 26808 2826 26817 2833
rect 26817 2826 26851 2833
rect 26851 2826 26860 2833
rect 26808 2788 26860 2826
rect 26808 2781 26817 2788
rect 26817 2781 26851 2788
rect 26851 2781 26860 2788
rect 27068 2826 27077 2833
rect 27077 2826 27111 2833
rect 27111 2826 27120 2833
rect 27068 2788 27120 2826
rect 27068 2781 27077 2788
rect 27077 2781 27111 2788
rect 27111 2781 27120 2788
rect 26678 2512 26730 2517
rect 26678 2478 26687 2512
rect 26687 2478 26721 2512
rect 26721 2478 26730 2512
rect 26678 2465 26730 2478
rect 26678 2440 26730 2453
rect 26678 2406 26687 2440
rect 26687 2406 26721 2440
rect 26721 2406 26730 2440
rect 26678 2401 26730 2406
rect 26808 2512 26860 2517
rect 26808 2478 26817 2512
rect 26817 2478 26851 2512
rect 26851 2478 26860 2512
rect 26808 2465 26860 2478
rect 26808 2440 26860 2453
rect 26808 2406 26817 2440
rect 26817 2406 26851 2440
rect 26851 2406 26860 2440
rect 26808 2401 26860 2406
rect 12596 2266 12648 2318
rect 24188 2266 24240 2318
rect 12897 2109 12949 2161
rect 13266 2109 13318 2161
rect 13656 2109 13708 2161
rect 14046 2109 14098 2161
rect 14436 2109 14488 2161
rect 14826 2109 14878 2161
rect 15216 2109 15268 2161
rect 15671 2109 15723 2161
rect 24489 2109 24541 2161
rect 24858 2109 24910 2161
rect 25248 2109 25300 2161
rect 25638 2109 25690 2161
rect 26028 2109 26080 2161
rect 26418 2109 26470 2161
rect 26808 2109 26860 2161
rect 27263 2109 27315 2161
rect 13266 1838 13275 1865
rect 13275 1838 13309 1865
rect 13309 1838 13318 1865
rect 13266 1813 13318 1838
rect 13266 1800 13318 1801
rect 13266 1766 13275 1800
rect 13275 1766 13309 1800
rect 13309 1766 13318 1800
rect 13266 1749 13318 1766
rect 13266 1728 13318 1737
rect 13266 1694 13275 1728
rect 13275 1694 13309 1728
rect 13309 1694 13318 1728
rect 13266 1685 13318 1694
rect 13266 1656 13318 1673
rect 13266 1622 13275 1656
rect 13275 1622 13309 1656
rect 13309 1622 13318 1656
rect 13266 1621 13318 1622
rect 13266 1584 13318 1609
rect 13266 1557 13275 1584
rect 13275 1557 13309 1584
rect 13309 1557 13318 1584
rect 13656 1838 13665 1865
rect 13665 1838 13699 1865
rect 13699 1838 13708 1865
rect 13656 1813 13708 1838
rect 13656 1800 13708 1801
rect 13656 1766 13665 1800
rect 13665 1766 13699 1800
rect 13699 1766 13708 1800
rect 13656 1749 13708 1766
rect 13656 1728 13708 1737
rect 13656 1694 13665 1728
rect 13665 1694 13699 1728
rect 13699 1694 13708 1728
rect 13656 1685 13708 1694
rect 13656 1656 13708 1673
rect 13656 1622 13665 1656
rect 13665 1622 13699 1656
rect 13699 1622 13708 1656
rect 13656 1621 13708 1622
rect 13656 1584 13708 1609
rect 13656 1557 13665 1584
rect 13665 1557 13699 1584
rect 13699 1557 13708 1584
rect 13136 1180 13188 1189
rect 13136 1146 13145 1180
rect 13145 1146 13179 1180
rect 13179 1146 13188 1180
rect 13136 1137 13188 1146
rect 13266 1180 13318 1189
rect 13266 1146 13275 1180
rect 13275 1146 13309 1180
rect 13309 1146 13318 1180
rect 13266 1137 13318 1146
rect 14046 1838 14055 1865
rect 14055 1838 14089 1865
rect 14089 1838 14098 1865
rect 14046 1813 14098 1838
rect 14046 1800 14098 1801
rect 14046 1766 14055 1800
rect 14055 1766 14089 1800
rect 14089 1766 14098 1800
rect 14046 1749 14098 1766
rect 14046 1728 14098 1737
rect 14046 1694 14055 1728
rect 14055 1694 14089 1728
rect 14089 1694 14098 1728
rect 14046 1685 14098 1694
rect 14046 1656 14098 1673
rect 14046 1622 14055 1656
rect 14055 1622 14089 1656
rect 14089 1622 14098 1656
rect 14046 1621 14098 1622
rect 14046 1584 14098 1609
rect 14046 1557 14055 1584
rect 14055 1557 14089 1584
rect 14089 1557 14098 1584
rect 13526 1180 13578 1189
rect 13526 1146 13535 1180
rect 13535 1146 13569 1180
rect 13569 1146 13578 1180
rect 13526 1137 13578 1146
rect 13656 1180 13708 1189
rect 13656 1146 13665 1180
rect 13665 1146 13699 1180
rect 13699 1146 13708 1180
rect 13656 1137 13708 1146
rect 14436 1838 14445 1865
rect 14445 1838 14479 1865
rect 14479 1838 14488 1865
rect 14436 1813 14488 1838
rect 14436 1800 14488 1801
rect 14436 1766 14445 1800
rect 14445 1766 14479 1800
rect 14479 1766 14488 1800
rect 14436 1749 14488 1766
rect 14436 1728 14488 1737
rect 14436 1694 14445 1728
rect 14445 1694 14479 1728
rect 14479 1694 14488 1728
rect 14436 1685 14488 1694
rect 14436 1656 14488 1673
rect 14436 1622 14445 1656
rect 14445 1622 14479 1656
rect 14479 1622 14488 1656
rect 14436 1621 14488 1622
rect 14436 1584 14488 1609
rect 14436 1557 14445 1584
rect 14445 1557 14479 1584
rect 14479 1557 14488 1584
rect 13916 1180 13968 1189
rect 13916 1146 13925 1180
rect 13925 1146 13959 1180
rect 13959 1146 13968 1180
rect 13916 1137 13968 1146
rect 14046 1180 14098 1189
rect 14046 1146 14055 1180
rect 14055 1146 14089 1180
rect 14089 1146 14098 1180
rect 14046 1137 14098 1146
rect 14826 1838 14835 1865
rect 14835 1838 14869 1865
rect 14869 1838 14878 1865
rect 14826 1813 14878 1838
rect 14826 1800 14878 1801
rect 14826 1766 14835 1800
rect 14835 1766 14869 1800
rect 14869 1766 14878 1800
rect 14826 1749 14878 1766
rect 14826 1728 14878 1737
rect 14826 1694 14835 1728
rect 14835 1694 14869 1728
rect 14869 1694 14878 1728
rect 14826 1685 14878 1694
rect 14826 1656 14878 1673
rect 14826 1622 14835 1656
rect 14835 1622 14869 1656
rect 14869 1622 14878 1656
rect 14826 1621 14878 1622
rect 14826 1584 14878 1609
rect 14826 1557 14835 1584
rect 14835 1557 14869 1584
rect 14869 1557 14878 1584
rect 14306 1180 14358 1189
rect 14306 1146 14315 1180
rect 14315 1146 14349 1180
rect 14349 1146 14358 1180
rect 14306 1137 14358 1146
rect 14436 1180 14488 1189
rect 14436 1146 14445 1180
rect 14445 1146 14479 1180
rect 14479 1146 14488 1180
rect 14436 1137 14488 1146
rect 15216 1838 15225 1865
rect 15225 1838 15259 1865
rect 15259 1838 15268 1865
rect 15216 1813 15268 1838
rect 15216 1800 15268 1801
rect 15216 1766 15225 1800
rect 15225 1766 15259 1800
rect 15259 1766 15268 1800
rect 15216 1749 15268 1766
rect 15216 1728 15268 1737
rect 15216 1694 15225 1728
rect 15225 1694 15259 1728
rect 15259 1694 15268 1728
rect 15216 1685 15268 1694
rect 15216 1656 15268 1673
rect 15216 1622 15225 1656
rect 15225 1622 15259 1656
rect 15259 1622 15268 1656
rect 15216 1621 15268 1622
rect 15216 1584 15268 1609
rect 15216 1557 15225 1584
rect 15225 1557 15259 1584
rect 15259 1557 15268 1584
rect 14696 1180 14748 1189
rect 14696 1146 14705 1180
rect 14705 1146 14739 1180
rect 14739 1146 14748 1180
rect 14696 1137 14748 1146
rect 14826 1180 14878 1189
rect 14826 1146 14835 1180
rect 14835 1146 14869 1180
rect 14869 1146 14878 1180
rect 14826 1137 14878 1146
rect 24858 1838 24867 1865
rect 24867 1838 24901 1865
rect 24901 1838 24910 1865
rect 24858 1813 24910 1838
rect 24858 1800 24910 1801
rect 24858 1766 24867 1800
rect 24867 1766 24901 1800
rect 24901 1766 24910 1800
rect 24858 1749 24910 1766
rect 24858 1728 24910 1737
rect 24858 1694 24867 1728
rect 24867 1694 24901 1728
rect 24901 1694 24910 1728
rect 24858 1685 24910 1694
rect 24858 1656 24910 1673
rect 24858 1622 24867 1656
rect 24867 1622 24901 1656
rect 24901 1622 24910 1656
rect 24858 1621 24910 1622
rect 24858 1584 24910 1609
rect 24858 1557 24867 1584
rect 24867 1557 24901 1584
rect 24901 1557 24910 1584
rect 15086 1180 15138 1189
rect 15086 1146 15095 1180
rect 15095 1146 15129 1180
rect 15129 1146 15138 1180
rect 15086 1137 15138 1146
rect 15216 1180 15268 1189
rect 15216 1146 15225 1180
rect 15225 1146 15259 1180
rect 15259 1146 15268 1180
rect 15216 1137 15268 1146
rect 25248 1838 25257 1865
rect 25257 1838 25291 1865
rect 25291 1838 25300 1865
rect 25248 1813 25300 1838
rect 25248 1800 25300 1801
rect 25248 1766 25257 1800
rect 25257 1766 25291 1800
rect 25291 1766 25300 1800
rect 25248 1749 25300 1766
rect 25248 1728 25300 1737
rect 25248 1694 25257 1728
rect 25257 1694 25291 1728
rect 25291 1694 25300 1728
rect 25248 1685 25300 1694
rect 25248 1656 25300 1673
rect 25248 1622 25257 1656
rect 25257 1622 25291 1656
rect 25291 1622 25300 1656
rect 25248 1621 25300 1622
rect 25248 1584 25300 1609
rect 25248 1557 25257 1584
rect 25257 1557 25291 1584
rect 25291 1557 25300 1584
rect 15476 1180 15528 1189
rect 15476 1146 15485 1180
rect 15485 1146 15519 1180
rect 15519 1146 15528 1180
rect 15476 1137 15528 1146
rect 24728 1180 24780 1189
rect 24728 1146 24737 1180
rect 24737 1146 24771 1180
rect 24771 1146 24780 1180
rect 24728 1137 24780 1146
rect 24858 1180 24910 1189
rect 24858 1146 24867 1180
rect 24867 1146 24901 1180
rect 24901 1146 24910 1180
rect 24858 1137 24910 1146
rect 25638 1838 25647 1865
rect 25647 1838 25681 1865
rect 25681 1838 25690 1865
rect 25638 1813 25690 1838
rect 25638 1800 25690 1801
rect 25638 1766 25647 1800
rect 25647 1766 25681 1800
rect 25681 1766 25690 1800
rect 25638 1749 25690 1766
rect 25638 1728 25690 1737
rect 25638 1694 25647 1728
rect 25647 1694 25681 1728
rect 25681 1694 25690 1728
rect 25638 1685 25690 1694
rect 25638 1656 25690 1673
rect 25638 1622 25647 1656
rect 25647 1622 25681 1656
rect 25681 1622 25690 1656
rect 25638 1621 25690 1622
rect 25638 1584 25690 1609
rect 25638 1557 25647 1584
rect 25647 1557 25681 1584
rect 25681 1557 25690 1584
rect 25118 1180 25170 1189
rect 25118 1146 25127 1180
rect 25127 1146 25161 1180
rect 25161 1146 25170 1180
rect 25118 1137 25170 1146
rect 25248 1180 25300 1189
rect 25248 1146 25257 1180
rect 25257 1146 25291 1180
rect 25291 1146 25300 1180
rect 25248 1137 25300 1146
rect 26028 1838 26037 1865
rect 26037 1838 26071 1865
rect 26071 1838 26080 1865
rect 26028 1813 26080 1838
rect 26028 1800 26080 1801
rect 26028 1766 26037 1800
rect 26037 1766 26071 1800
rect 26071 1766 26080 1800
rect 26028 1749 26080 1766
rect 26028 1728 26080 1737
rect 26028 1694 26037 1728
rect 26037 1694 26071 1728
rect 26071 1694 26080 1728
rect 26028 1685 26080 1694
rect 26028 1656 26080 1673
rect 26028 1622 26037 1656
rect 26037 1622 26071 1656
rect 26071 1622 26080 1656
rect 26028 1621 26080 1622
rect 26028 1584 26080 1609
rect 26028 1557 26037 1584
rect 26037 1557 26071 1584
rect 26071 1557 26080 1584
rect 25508 1180 25560 1189
rect 25508 1146 25517 1180
rect 25517 1146 25551 1180
rect 25551 1146 25560 1180
rect 25508 1137 25560 1146
rect 25638 1180 25690 1189
rect 25638 1146 25647 1180
rect 25647 1146 25681 1180
rect 25681 1146 25690 1180
rect 25638 1137 25690 1146
rect 26418 1838 26427 1865
rect 26427 1838 26461 1865
rect 26461 1838 26470 1865
rect 26418 1813 26470 1838
rect 26418 1800 26470 1801
rect 26418 1766 26427 1800
rect 26427 1766 26461 1800
rect 26461 1766 26470 1800
rect 26418 1749 26470 1766
rect 26418 1728 26470 1737
rect 26418 1694 26427 1728
rect 26427 1694 26461 1728
rect 26461 1694 26470 1728
rect 26418 1685 26470 1694
rect 26418 1656 26470 1673
rect 26418 1622 26427 1656
rect 26427 1622 26461 1656
rect 26461 1622 26470 1656
rect 26418 1621 26470 1622
rect 26418 1584 26470 1609
rect 26418 1557 26427 1584
rect 26427 1557 26461 1584
rect 26461 1557 26470 1584
rect 25898 1180 25950 1189
rect 25898 1146 25907 1180
rect 25907 1146 25941 1180
rect 25941 1146 25950 1180
rect 25898 1137 25950 1146
rect 26028 1180 26080 1189
rect 26028 1146 26037 1180
rect 26037 1146 26071 1180
rect 26071 1146 26080 1180
rect 26028 1137 26080 1146
rect 26808 1838 26817 1865
rect 26817 1838 26851 1865
rect 26851 1838 26860 1865
rect 26808 1813 26860 1838
rect 26808 1800 26860 1801
rect 26808 1766 26817 1800
rect 26817 1766 26851 1800
rect 26851 1766 26860 1800
rect 26808 1749 26860 1766
rect 26808 1728 26860 1737
rect 26808 1694 26817 1728
rect 26817 1694 26851 1728
rect 26851 1694 26860 1728
rect 26808 1685 26860 1694
rect 26808 1656 26860 1673
rect 26808 1622 26817 1656
rect 26817 1622 26851 1656
rect 26851 1622 26860 1656
rect 26808 1621 26860 1622
rect 26808 1584 26860 1609
rect 26808 1557 26817 1584
rect 26817 1557 26851 1584
rect 26851 1557 26860 1584
rect 26288 1180 26340 1189
rect 26288 1146 26297 1180
rect 26297 1146 26331 1180
rect 26331 1146 26340 1180
rect 26288 1137 26340 1146
rect 26418 1180 26470 1189
rect 26418 1146 26427 1180
rect 26427 1146 26461 1180
rect 26461 1146 26470 1180
rect 26418 1137 26470 1146
rect 26678 1180 26730 1189
rect 26678 1146 26687 1180
rect 26687 1146 26721 1180
rect 26721 1146 26730 1180
rect 26678 1137 26730 1146
rect 26808 1180 26860 1189
rect 26808 1146 26817 1180
rect 26817 1146 26851 1180
rect 26851 1146 26860 1180
rect 26808 1137 26860 1146
rect 27068 1180 27120 1189
rect 27068 1146 27077 1180
rect 27077 1146 27111 1180
rect 27111 1146 27120 1180
rect 27068 1137 27120 1146
rect 12504 864 12556 916
rect 13331 907 13383 916
rect 13331 873 13340 907
rect 13340 873 13374 907
rect 13374 873 13383 907
rect 13331 864 13383 873
rect 13721 907 13773 916
rect 13721 873 13730 907
rect 13730 873 13764 907
rect 13764 873 13773 907
rect 13721 864 13773 873
rect 14111 907 14163 916
rect 14111 873 14120 907
rect 14120 873 14154 907
rect 14154 873 14163 907
rect 14111 864 14163 873
rect 14501 907 14553 916
rect 14501 873 14510 907
rect 14510 873 14544 907
rect 14544 873 14553 907
rect 14501 864 14553 873
rect 14891 907 14943 916
rect 14891 873 14900 907
rect 14900 873 14934 907
rect 14934 873 14943 907
rect 14891 864 14943 873
rect 15281 907 15333 916
rect 15281 873 15290 907
rect 15290 873 15324 907
rect 15324 873 15333 907
rect 15281 864 15333 873
rect 24096 864 24148 916
rect 24923 907 24975 916
rect 24923 873 24932 907
rect 24932 873 24966 907
rect 24966 873 24975 907
rect 24923 864 24975 873
rect 25313 907 25365 916
rect 25313 873 25322 907
rect 25322 873 25356 907
rect 25356 873 25365 907
rect 25313 864 25365 873
rect 25703 907 25755 916
rect 25703 873 25712 907
rect 25712 873 25746 907
rect 25746 873 25755 907
rect 25703 864 25755 873
rect 26093 907 26145 916
rect 26093 873 26102 907
rect 26102 873 26136 907
rect 26136 873 26145 907
rect 26093 864 26145 873
rect 26483 907 26535 916
rect 26483 873 26492 907
rect 26492 873 26526 907
rect 26526 873 26535 907
rect 26483 864 26535 873
rect 26873 907 26925 916
rect 26873 873 26882 907
rect 26882 873 26916 907
rect 26916 873 26925 907
rect 26873 864 26925 873
rect 12833 731 12885 783
rect 12897 731 12949 783
rect 12961 731 13013 783
rect 13657 774 13709 783
rect 13657 740 13658 774
rect 13658 740 13692 774
rect 13692 740 13709 774
rect 13657 731 13709 740
rect 13721 774 13773 783
rect 13721 740 13730 774
rect 13730 740 13764 774
rect 13764 740 13773 774
rect 13721 731 13773 740
rect 13785 774 13837 783
rect 14437 774 14489 783
rect 13785 740 13802 774
rect 13802 740 13836 774
rect 13836 740 13837 774
rect 14437 740 14438 774
rect 14438 740 14472 774
rect 14472 740 14489 774
rect 13785 731 13837 740
rect 14437 731 14489 740
rect 14501 774 14553 783
rect 14501 740 14510 774
rect 14510 740 14544 774
rect 14544 740 14553 774
rect 14501 731 14553 740
rect 14565 774 14617 783
rect 15217 774 15269 783
rect 14565 740 14582 774
rect 14582 740 14616 774
rect 14616 740 14617 774
rect 15217 740 15218 774
rect 15218 740 15252 774
rect 15252 740 15269 774
rect 14565 731 14617 740
rect 15217 731 15269 740
rect 15281 774 15333 783
rect 15281 740 15290 774
rect 15290 740 15324 774
rect 15324 740 15333 774
rect 15281 731 15333 740
rect 15345 774 15397 783
rect 15345 740 15362 774
rect 15362 740 15396 774
rect 15396 740 15397 774
rect 15345 731 15397 740
rect 24425 731 24477 783
rect 24489 731 24541 783
rect 24553 731 24605 783
rect 25249 774 25301 783
rect 25249 740 25250 774
rect 25250 740 25284 774
rect 25284 740 25301 774
rect 25249 731 25301 740
rect 25313 774 25365 783
rect 25313 740 25322 774
rect 25322 740 25356 774
rect 25356 740 25365 774
rect 25313 731 25365 740
rect 25377 774 25429 783
rect 26029 774 26081 783
rect 25377 740 25394 774
rect 25394 740 25428 774
rect 25428 740 25429 774
rect 26029 740 26030 774
rect 26030 740 26064 774
rect 26064 740 26081 774
rect 25377 731 25429 740
rect 26029 731 26081 740
rect 26093 774 26145 783
rect 26093 740 26102 774
rect 26102 740 26136 774
rect 26136 740 26145 774
rect 26093 731 26145 740
rect 26157 774 26209 783
rect 26809 774 26861 783
rect 26157 740 26174 774
rect 26174 740 26208 774
rect 26208 740 26209 774
rect 26809 740 26810 774
rect 26810 740 26844 774
rect 26844 740 26861 774
rect 26157 731 26209 740
rect 26809 731 26861 740
rect 26873 774 26925 783
rect 26873 740 26882 774
rect 26882 740 26916 774
rect 26916 740 26925 774
rect 26873 731 26925 740
rect 26937 774 26989 783
rect 26937 740 26954 774
rect 26954 740 26988 774
rect 26988 740 26989 774
rect 26937 731 26989 740
<< metal2 >>
rect 12823 5497 13023 5509
rect 12823 5495 12855 5497
rect 12911 5495 12935 5497
rect 12991 5495 13023 5497
rect 12823 5443 12833 5495
rect 13013 5443 13023 5495
rect 12823 5441 12855 5443
rect 12911 5441 12935 5443
rect 12991 5441 13023 5443
rect 12823 5429 13023 5441
rect 13647 5497 13847 5509
rect 13647 5495 13679 5497
rect 13735 5495 13759 5497
rect 13815 5495 13847 5497
rect 13647 5443 13657 5495
rect 13837 5443 13847 5495
rect 13647 5441 13679 5443
rect 13735 5441 13759 5443
rect 13815 5441 13847 5443
rect 13647 5429 13847 5441
rect 14427 5497 14627 5509
rect 14427 5495 14459 5497
rect 14515 5495 14539 5497
rect 14595 5495 14627 5497
rect 14427 5443 14437 5495
rect 14617 5443 14627 5495
rect 14427 5441 14459 5443
rect 14515 5441 14539 5443
rect 14595 5441 14627 5443
rect 14427 5429 14627 5441
rect 15207 5497 15407 5509
rect 15207 5495 15239 5497
rect 15295 5495 15319 5497
rect 15375 5495 15407 5497
rect 15207 5443 15217 5495
rect 15397 5443 15407 5495
rect 15207 5441 15239 5443
rect 15295 5441 15319 5443
rect 15375 5441 15407 5443
rect 15207 5429 15407 5441
rect 24415 5497 24615 5509
rect 24415 5495 24447 5497
rect 24503 5495 24527 5497
rect 24583 5495 24615 5497
rect 24415 5443 24425 5495
rect 24605 5443 24615 5495
rect 24415 5441 24447 5443
rect 24503 5441 24527 5443
rect 24583 5441 24615 5443
rect 24415 5429 24615 5441
rect 25239 5497 25439 5509
rect 25239 5495 25271 5497
rect 25327 5495 25351 5497
rect 25407 5495 25439 5497
rect 25239 5443 25249 5495
rect 25429 5443 25439 5495
rect 25239 5441 25271 5443
rect 25327 5441 25351 5443
rect 25407 5441 25439 5443
rect 25239 5429 25439 5441
rect 26019 5497 26219 5509
rect 26019 5495 26051 5497
rect 26107 5495 26131 5497
rect 26187 5495 26219 5497
rect 26019 5443 26029 5495
rect 26209 5443 26219 5495
rect 26019 5441 26051 5443
rect 26107 5441 26131 5443
rect 26187 5441 26219 5443
rect 26019 5429 26219 5441
rect 26799 5497 26999 5509
rect 26799 5495 26831 5497
rect 26887 5495 26911 5497
rect 26967 5495 26999 5497
rect 26799 5443 26809 5495
rect 26989 5443 26999 5495
rect 26799 5441 26831 5443
rect 26887 5441 26911 5443
rect 26967 5441 26999 5443
rect 26799 5429 26999 5441
rect 12493 5364 12567 5369
rect 12493 5308 12502 5364
rect 12558 5308 12567 5364
rect 12493 5303 12567 5308
rect 13000 5364 13134 5369
rect 13000 5362 13039 5364
rect 13095 5362 13134 5364
rect 13000 5310 13009 5362
rect 13125 5310 13134 5362
rect 13000 5308 13039 5310
rect 13095 5308 13134 5310
rect 13000 5303 13134 5308
rect 13320 5364 13394 5369
rect 13320 5308 13329 5364
rect 13385 5308 13394 5364
rect 13320 5303 13394 5308
rect 13710 5364 13784 5369
rect 13710 5308 13719 5364
rect 13775 5308 13784 5364
rect 13710 5303 13784 5308
rect 14100 5364 14174 5369
rect 14100 5308 14109 5364
rect 14165 5308 14174 5364
rect 14100 5303 14174 5308
rect 14490 5364 14564 5369
rect 14490 5308 14499 5364
rect 14555 5308 14564 5364
rect 14490 5303 14564 5308
rect 14880 5364 14954 5369
rect 14880 5308 14889 5364
rect 14945 5308 14954 5364
rect 14880 5303 14954 5308
rect 24085 5364 24159 5369
rect 24085 5308 24094 5364
rect 24150 5308 24159 5364
rect 24085 5303 24159 5308
rect 24592 5364 24726 5369
rect 24592 5362 24631 5364
rect 24687 5362 24726 5364
rect 24592 5310 24601 5362
rect 24717 5310 24726 5362
rect 24592 5308 24631 5310
rect 24687 5308 24726 5310
rect 24592 5303 24726 5308
rect 24912 5364 24986 5369
rect 24912 5308 24921 5364
rect 24977 5308 24986 5364
rect 24912 5303 24986 5308
rect 25302 5364 25376 5369
rect 25302 5308 25311 5364
rect 25367 5308 25376 5364
rect 25302 5303 25376 5308
rect 25692 5364 25766 5369
rect 25692 5308 25701 5364
rect 25757 5308 25766 5364
rect 25692 5303 25766 5308
rect 26082 5364 26156 5369
rect 26082 5308 26091 5364
rect 26147 5308 26156 5364
rect 26082 5303 26156 5308
rect 26472 5364 26546 5369
rect 26472 5308 26481 5364
rect 26537 5308 26546 5364
rect 26472 5303 26546 5308
rect 12503 923 12557 5303
rect 13000 5217 13064 5303
rect 13000 5165 13006 5217
rect 13058 5165 13064 5217
rect 13000 5153 13064 5165
rect 13000 5101 13006 5153
rect 13058 5101 13064 5153
rect 13000 5089 13064 5101
rect 13000 5037 13006 5089
rect 13058 5037 13064 5089
rect 13000 5025 13064 5037
rect 13000 4973 13006 5025
rect 13058 4973 13064 5025
rect 13125 5091 13199 5113
rect 13125 5035 13134 5091
rect 13190 5035 13199 5091
rect 13125 5013 13199 5035
rect 13385 5091 13459 5113
rect 13385 5035 13394 5091
rect 13450 5035 13459 5091
rect 13385 5013 13459 5035
rect 13515 5091 13589 5113
rect 13515 5035 13524 5091
rect 13580 5035 13589 5091
rect 13515 5013 13589 5035
rect 13775 5091 13849 5113
rect 13775 5035 13784 5091
rect 13840 5035 13849 5091
rect 13775 5013 13849 5035
rect 13905 5091 13979 5113
rect 13905 5035 13914 5091
rect 13970 5035 13979 5091
rect 13905 5013 13979 5035
rect 14165 5091 14239 5113
rect 14165 5035 14174 5091
rect 14230 5035 14239 5091
rect 14165 5013 14239 5035
rect 14295 5091 14369 5113
rect 14295 5035 14304 5091
rect 14360 5035 14369 5091
rect 14295 5013 14369 5035
rect 14555 5091 14629 5113
rect 14555 5035 14564 5091
rect 14620 5035 14629 5091
rect 14555 5013 14629 5035
rect 14685 5091 14759 5113
rect 14685 5035 14694 5091
rect 14750 5035 14759 5091
rect 14685 5013 14759 5035
rect 14945 5091 15019 5113
rect 14945 5035 14954 5091
rect 15010 5035 15019 5091
rect 14945 5013 15019 5035
rect 15075 5091 15149 5113
rect 15075 5035 15084 5091
rect 15140 5035 15149 5091
rect 15075 5013 15149 5035
rect 13000 4961 13064 4973
rect 13000 4909 13006 4961
rect 13058 4909 13064 4961
rect 12891 4117 12955 4123
rect 12891 4065 12897 4117
rect 12949 4065 12955 4117
rect 12590 3960 12654 3961
rect 12590 3908 12596 3960
rect 12648 3908 12654 3960
rect 12590 3907 12654 3908
rect 12595 3405 12649 3907
rect 12585 3400 12659 3405
rect 12585 3344 12594 3400
rect 12650 3344 12659 3400
rect 12585 3339 12659 3344
rect 12595 2319 12649 3339
rect 12677 3274 12751 3279
rect 12677 3218 12686 3274
rect 12742 3218 12751 3274
rect 12677 3213 12751 3218
rect 12687 3013 12741 3213
rect 12677 3008 12751 3013
rect 12677 2952 12686 3008
rect 12742 2952 12751 3008
rect 12677 2947 12751 2952
rect 12590 2318 12654 2319
rect 12590 2266 12596 2318
rect 12648 2266 12654 2318
rect 12590 2265 12654 2266
rect 12891 2161 12955 4065
rect 13000 3477 13064 4909
rect 15207 4926 15407 4931
rect 15207 4870 15239 4926
rect 15295 4924 15319 4926
rect 15375 4925 15407 4926
rect 15375 4924 15518 4925
rect 15295 4872 15317 4924
rect 15375 4872 15381 4924
rect 15433 4872 15445 4924
rect 15497 4872 15518 4924
rect 15295 4870 15319 4872
rect 15375 4871 15518 4872
rect 15375 4870 15407 4871
rect 15207 4865 15407 4870
rect 15198 4781 15204 4833
rect 15256 4781 15262 4833
rect 13390 4669 13454 4688
rect 13390 4617 13396 4669
rect 13448 4617 13454 4669
rect 13390 4605 13454 4617
rect 13390 4553 13396 4605
rect 13448 4553 13454 4605
rect 13390 4541 13454 4553
rect 13390 4489 13396 4541
rect 13448 4489 13454 4541
rect 13390 4477 13454 4489
rect 13390 4425 13396 4477
rect 13448 4425 13454 4477
rect 13390 4413 13454 4425
rect 13390 4361 13396 4413
rect 13448 4361 13454 4413
rect 13390 4342 13454 4361
rect 13780 4669 13844 4688
rect 13780 4617 13786 4669
rect 13838 4617 13844 4669
rect 13780 4605 13844 4617
rect 13780 4553 13786 4605
rect 13838 4553 13844 4605
rect 13780 4541 13844 4553
rect 13780 4489 13786 4541
rect 13838 4489 13844 4541
rect 13780 4477 13844 4489
rect 13780 4425 13786 4477
rect 13838 4425 13844 4477
rect 13780 4413 13844 4425
rect 13780 4361 13786 4413
rect 13838 4361 13844 4413
rect 13780 4342 13844 4361
rect 14170 4669 14234 4688
rect 14170 4617 14176 4669
rect 14228 4617 14234 4669
rect 14170 4605 14234 4617
rect 14170 4553 14176 4605
rect 14228 4553 14234 4605
rect 14170 4541 14234 4553
rect 14170 4489 14176 4541
rect 14228 4489 14234 4541
rect 14170 4477 14234 4489
rect 14170 4425 14176 4477
rect 14228 4425 14234 4477
rect 14170 4413 14234 4425
rect 14170 4361 14176 4413
rect 14228 4361 14234 4413
rect 14170 4342 14234 4361
rect 14560 4669 14624 4688
rect 14560 4617 14566 4669
rect 14618 4617 14624 4669
rect 14560 4605 14624 4617
rect 14560 4553 14566 4605
rect 14618 4553 14624 4605
rect 14560 4541 14624 4553
rect 14560 4489 14566 4541
rect 14618 4489 14624 4541
rect 14560 4477 14624 4489
rect 14560 4425 14566 4477
rect 14618 4425 14624 4477
rect 14560 4413 14624 4425
rect 14560 4361 14566 4413
rect 14618 4361 14624 4413
rect 14560 4342 14624 4361
rect 14950 4669 15014 4688
rect 14950 4617 14956 4669
rect 15008 4617 15014 4669
rect 14950 4605 15014 4617
rect 14950 4553 14956 4605
rect 15008 4553 15014 4605
rect 14950 4541 15014 4553
rect 14950 4489 14956 4541
rect 15008 4489 15014 4541
rect 14950 4477 15014 4489
rect 14950 4425 14956 4477
rect 15008 4425 15014 4477
rect 14950 4413 15014 4425
rect 14950 4361 14956 4413
rect 15008 4361 15014 4413
rect 15205 4397 15245 4781
rect 15298 4685 15338 4865
rect 15475 4685 15515 4871
rect 15284 4633 15290 4685
rect 15342 4633 15348 4685
rect 15464 4633 15470 4685
rect 15522 4633 15528 4685
rect 14950 4342 15014 4361
rect 15194 4345 15200 4397
rect 15252 4345 15258 4397
rect 15373 4391 15439 4392
rect 13399 4123 13445 4342
rect 13789 4123 13835 4342
rect 14179 4123 14225 4342
rect 14569 4123 14615 4342
rect 14959 4123 15005 4342
rect 13390 4117 13454 4123
rect 13390 4065 13396 4117
rect 13448 4065 13454 4117
rect 13390 4059 13454 4065
rect 13780 4117 13844 4123
rect 13780 4065 13786 4117
rect 13838 4065 13844 4117
rect 13780 4059 13844 4065
rect 14170 4117 14234 4123
rect 14170 4065 14176 4117
rect 14228 4065 14234 4117
rect 14170 4059 14234 4065
rect 14560 4117 14624 4123
rect 14560 4065 14566 4117
rect 14618 4065 14624 4117
rect 14560 4059 14624 4065
rect 14950 4117 15014 4123
rect 14950 4065 14956 4117
rect 15008 4065 15014 4117
rect 14950 4059 15014 4065
rect 13399 3832 13445 4059
rect 13789 3832 13835 4059
rect 14179 3832 14225 4059
rect 14569 3832 14615 4059
rect 14959 3832 15005 4059
rect 13390 3825 13454 3832
rect 13390 3773 13396 3825
rect 13448 3773 13454 3825
rect 13390 3761 13454 3773
rect 13390 3709 13396 3761
rect 13448 3709 13454 3761
rect 13390 3702 13454 3709
rect 13520 3825 13584 3832
rect 13520 3773 13526 3825
rect 13578 3773 13584 3825
rect 13520 3761 13584 3773
rect 13520 3709 13526 3761
rect 13578 3709 13584 3761
rect 13520 3702 13584 3709
rect 13780 3825 13844 3832
rect 13780 3773 13786 3825
rect 13838 3773 13844 3825
rect 13780 3761 13844 3773
rect 13780 3709 13786 3761
rect 13838 3709 13844 3761
rect 13780 3702 13844 3709
rect 13910 3825 13974 3832
rect 13910 3773 13916 3825
rect 13968 3773 13974 3825
rect 13910 3761 13974 3773
rect 13910 3709 13916 3761
rect 13968 3709 13974 3761
rect 13910 3702 13974 3709
rect 14170 3825 14234 3832
rect 14170 3773 14176 3825
rect 14228 3773 14234 3825
rect 14170 3761 14234 3773
rect 14170 3709 14176 3761
rect 14228 3709 14234 3761
rect 14170 3702 14234 3709
rect 14300 3825 14364 3832
rect 14300 3773 14306 3825
rect 14358 3773 14364 3825
rect 14300 3761 14364 3773
rect 14300 3709 14306 3761
rect 14358 3709 14364 3761
rect 14300 3702 14364 3709
rect 14560 3825 14624 3832
rect 14560 3773 14566 3825
rect 14618 3773 14624 3825
rect 14560 3761 14624 3773
rect 14560 3709 14566 3761
rect 14618 3709 14624 3761
rect 14560 3702 14624 3709
rect 14690 3825 14754 3832
rect 14690 3773 14696 3825
rect 14748 3773 14754 3825
rect 14690 3761 14754 3773
rect 14690 3709 14696 3761
rect 14748 3709 14754 3761
rect 14690 3702 14754 3709
rect 14950 3825 15014 3832
rect 14950 3773 14956 3825
rect 15008 3773 15014 3825
rect 14950 3761 15014 3773
rect 14950 3709 14956 3761
rect 15008 3709 15014 3761
rect 14950 3702 15014 3709
rect 15080 3825 15144 3832
rect 15205 3829 15245 4345
rect 15373 4339 15380 4391
rect 15432 4339 15439 4391
rect 15373 4338 15439 4339
rect 15553 4391 15619 4392
rect 15553 4339 15560 4391
rect 15612 4339 15619 4391
rect 15553 4338 15619 4339
rect 15386 4296 15426 4338
rect 15566 4296 15606 4338
rect 15797 4297 15957 4302
rect 15373 4295 15439 4296
rect 15373 4243 15380 4295
rect 15432 4243 15439 4295
rect 15373 4242 15439 4243
rect 15553 4295 15619 4296
rect 15553 4243 15560 4295
rect 15612 4243 15619 4295
rect 15553 4242 15619 4243
rect 15386 3829 15426 4242
rect 15566 3829 15606 4242
rect 15797 4241 15809 4297
rect 15865 4295 15889 4297
rect 15871 4243 15883 4295
rect 15865 4241 15889 4243
rect 15945 4241 15957 4297
rect 15797 4236 15957 4241
rect 15665 4117 15729 4123
rect 15665 4065 15671 4117
rect 15723 4065 15729 4117
rect 15080 3773 15086 3825
rect 15138 3773 15144 3825
rect 15194 3777 15200 3829
rect 15252 3777 15258 3829
rect 15374 3777 15380 3829
rect 15432 3777 15438 3829
rect 15554 3777 15560 3829
rect 15612 3777 15618 3829
rect 15080 3761 15144 3773
rect 15080 3709 15086 3761
rect 15138 3709 15144 3761
rect 15080 3702 15144 3709
rect 15284 3705 15290 3757
rect 15342 3705 15348 3757
rect 15464 3705 15470 3757
rect 15522 3705 15528 3757
rect 13000 3425 13006 3477
rect 13058 3425 13064 3477
rect 13535 3469 13569 3702
rect 13925 3469 13959 3702
rect 14315 3469 14349 3702
rect 14705 3469 14739 3702
rect 15095 3469 15129 3702
rect 15294 3589 15334 3705
rect 15477 3595 15517 3705
rect 15467 3590 15637 3595
rect 15467 3589 15484 3590
rect 15294 3588 15484 3589
rect 15294 3536 15316 3588
rect 15368 3536 15380 3588
rect 15432 3536 15444 3588
rect 15294 3535 15484 3536
rect 15294 3533 15334 3535
rect 15467 3534 15484 3535
rect 15540 3534 15564 3590
rect 15620 3534 15637 3590
rect 15467 3529 15637 3534
rect 13000 3413 13064 3425
rect 13000 3361 13006 3413
rect 13058 3361 13064 3413
rect 13125 3447 13199 3469
rect 13125 3391 13134 3447
rect 13190 3391 13199 3447
rect 13125 3369 13199 3391
rect 13385 3447 13459 3469
rect 13385 3391 13394 3447
rect 13450 3391 13459 3447
rect 13385 3369 13459 3391
rect 13515 3447 13589 3469
rect 13515 3391 13524 3447
rect 13580 3391 13589 3447
rect 13515 3369 13589 3391
rect 13775 3447 13849 3469
rect 13775 3391 13784 3447
rect 13840 3391 13849 3447
rect 13775 3369 13849 3391
rect 13905 3447 13979 3469
rect 13905 3391 13914 3447
rect 13970 3391 13979 3447
rect 13905 3369 13979 3391
rect 14165 3447 14239 3469
rect 14165 3391 14174 3447
rect 14230 3391 14239 3447
rect 14165 3369 14239 3391
rect 14295 3447 14369 3469
rect 14295 3391 14304 3447
rect 14360 3391 14369 3447
rect 14295 3369 14369 3391
rect 14555 3447 14629 3469
rect 14555 3391 14564 3447
rect 14620 3391 14629 3447
rect 14555 3369 14629 3391
rect 14685 3447 14759 3469
rect 14685 3391 14694 3447
rect 14750 3391 14759 3447
rect 14685 3369 14759 3391
rect 14945 3447 15019 3469
rect 14945 3391 14954 3447
rect 15010 3391 15019 3447
rect 14945 3369 15019 3391
rect 15075 3447 15149 3469
rect 15075 3391 15084 3447
rect 15140 3391 15149 3447
rect 15075 3369 15149 3391
rect 13000 3354 13064 3361
rect 12992 3274 13066 3279
rect 12992 3218 13001 3274
rect 13057 3218 13066 3274
rect 12992 3213 13066 3218
rect 13320 3274 13394 3279
rect 13320 3218 13329 3274
rect 13385 3218 13394 3274
rect 13320 3213 13394 3218
rect 13710 3274 13784 3279
rect 13710 3218 13719 3274
rect 13775 3218 13784 3274
rect 13710 3213 13784 3218
rect 14100 3274 14174 3279
rect 14100 3218 14109 3274
rect 14165 3218 14174 3274
rect 14100 3213 14174 3218
rect 14490 3274 14564 3279
rect 14490 3218 14499 3274
rect 14555 3218 14564 3274
rect 14490 3213 14564 3218
rect 14880 3274 14954 3279
rect 14880 3218 14889 3274
rect 14945 3218 14954 3274
rect 14880 3213 14954 3218
rect 13257 3141 13457 3153
rect 13257 3139 13289 3141
rect 13345 3139 13369 3141
rect 13425 3139 13457 3141
rect 13257 3087 13267 3139
rect 13447 3087 13457 3139
rect 13257 3085 13289 3087
rect 13345 3085 13369 3087
rect 13425 3085 13457 3087
rect 13257 3073 13457 3085
rect 14037 3141 14237 3153
rect 14037 3139 14069 3141
rect 14125 3139 14149 3141
rect 14205 3139 14237 3141
rect 14037 3087 14047 3139
rect 14227 3087 14237 3139
rect 14037 3085 14069 3087
rect 14125 3085 14149 3087
rect 14205 3085 14237 3087
rect 14037 3073 14237 3085
rect 14817 3141 15017 3153
rect 14817 3139 14849 3141
rect 14905 3139 14929 3141
rect 14985 3139 15017 3141
rect 14817 3087 14827 3139
rect 15007 3087 15017 3139
rect 14817 3085 14849 3087
rect 14905 3085 14929 3087
rect 14985 3085 15017 3087
rect 14817 3073 15017 3085
rect 13320 3008 13394 3013
rect 13320 2952 13329 3008
rect 13385 2952 13394 3008
rect 13320 2947 13394 2952
rect 13710 3008 13784 3013
rect 13710 2952 13719 3008
rect 13775 2952 13784 3008
rect 13710 2947 13784 2952
rect 14100 3008 14174 3013
rect 14100 2952 14109 3008
rect 14165 2952 14174 3008
rect 14100 2947 14174 2952
rect 14490 3008 14564 3013
rect 14490 2952 14499 3008
rect 14555 2952 14564 3008
rect 14490 2947 14564 2952
rect 14880 3008 14954 3013
rect 14880 2952 14889 3008
rect 14945 2952 14954 3008
rect 14880 2947 14954 2952
rect 15270 3008 15344 3013
rect 15270 2952 15279 3008
rect 15335 2952 15344 3008
rect 15270 2947 15344 2952
rect 13125 2835 13199 2857
rect 13125 2779 13134 2835
rect 13190 2779 13199 2835
rect 13125 2757 13199 2779
rect 13255 2835 13329 2857
rect 13255 2779 13264 2835
rect 13320 2779 13329 2835
rect 13255 2757 13329 2779
rect 13515 2835 13589 2857
rect 13515 2779 13524 2835
rect 13580 2779 13589 2835
rect 13515 2757 13589 2779
rect 13645 2835 13719 2857
rect 13645 2779 13654 2835
rect 13710 2779 13719 2835
rect 13645 2757 13719 2779
rect 13905 2835 13979 2857
rect 13905 2779 13914 2835
rect 13970 2779 13979 2835
rect 13905 2757 13979 2779
rect 14035 2835 14109 2857
rect 14035 2779 14044 2835
rect 14100 2779 14109 2835
rect 14035 2757 14109 2779
rect 14295 2835 14369 2857
rect 14295 2779 14304 2835
rect 14360 2779 14369 2835
rect 14295 2757 14369 2779
rect 14425 2835 14499 2857
rect 14425 2779 14434 2835
rect 14490 2779 14499 2835
rect 14425 2757 14499 2779
rect 14685 2835 14759 2857
rect 14685 2779 14694 2835
rect 14750 2779 14759 2835
rect 14685 2757 14759 2779
rect 14815 2835 14889 2857
rect 14815 2779 14824 2835
rect 14880 2779 14889 2835
rect 14815 2757 14889 2779
rect 15075 2835 15149 2857
rect 15075 2779 15084 2835
rect 15140 2779 15149 2835
rect 15075 2757 15149 2779
rect 15205 2835 15279 2857
rect 15205 2779 15214 2835
rect 15270 2779 15279 2835
rect 15205 2757 15279 2779
rect 15465 2835 15539 2857
rect 15465 2779 15474 2835
rect 15530 2779 15539 2835
rect 15465 2757 15539 2779
rect 13145 2524 13179 2757
rect 13535 2524 13569 2757
rect 13925 2524 13959 2757
rect 14315 2524 14349 2757
rect 14705 2524 14739 2757
rect 15095 2524 15129 2757
rect 13130 2517 13194 2524
rect 13130 2465 13136 2517
rect 13188 2465 13194 2517
rect 13130 2453 13194 2465
rect 13130 2401 13136 2453
rect 13188 2401 13194 2453
rect 13130 2394 13194 2401
rect 13260 2517 13324 2524
rect 13260 2465 13266 2517
rect 13318 2465 13324 2517
rect 13260 2453 13324 2465
rect 13260 2401 13266 2453
rect 13318 2401 13324 2453
rect 13260 2394 13324 2401
rect 13520 2517 13584 2524
rect 13520 2465 13526 2517
rect 13578 2465 13584 2517
rect 13520 2453 13584 2465
rect 13520 2401 13526 2453
rect 13578 2401 13584 2453
rect 13520 2394 13584 2401
rect 13650 2517 13714 2524
rect 13650 2465 13656 2517
rect 13708 2465 13714 2517
rect 13650 2453 13714 2465
rect 13650 2401 13656 2453
rect 13708 2401 13714 2453
rect 13650 2394 13714 2401
rect 13910 2517 13974 2524
rect 13910 2465 13916 2517
rect 13968 2465 13974 2517
rect 13910 2453 13974 2465
rect 13910 2401 13916 2453
rect 13968 2401 13974 2453
rect 13910 2394 13974 2401
rect 14040 2517 14104 2524
rect 14040 2465 14046 2517
rect 14098 2465 14104 2517
rect 14040 2453 14104 2465
rect 14040 2401 14046 2453
rect 14098 2401 14104 2453
rect 14040 2394 14104 2401
rect 14300 2517 14364 2524
rect 14300 2465 14306 2517
rect 14358 2465 14364 2517
rect 14300 2453 14364 2465
rect 14300 2401 14306 2453
rect 14358 2401 14364 2453
rect 14300 2394 14364 2401
rect 14430 2517 14494 2524
rect 14430 2465 14436 2517
rect 14488 2465 14494 2517
rect 14430 2453 14494 2465
rect 14430 2401 14436 2453
rect 14488 2401 14494 2453
rect 14430 2394 14494 2401
rect 14690 2517 14754 2524
rect 14690 2465 14696 2517
rect 14748 2465 14754 2517
rect 14690 2453 14754 2465
rect 14690 2401 14696 2453
rect 14748 2401 14754 2453
rect 14690 2394 14754 2401
rect 14820 2517 14884 2524
rect 14820 2465 14826 2517
rect 14878 2465 14884 2517
rect 14820 2453 14884 2465
rect 14820 2401 14826 2453
rect 14878 2401 14884 2453
rect 14820 2394 14884 2401
rect 15080 2517 15144 2524
rect 15080 2465 15086 2517
rect 15138 2465 15144 2517
rect 15080 2453 15144 2465
rect 15080 2401 15086 2453
rect 15138 2401 15144 2453
rect 15080 2394 15144 2401
rect 15210 2517 15274 2524
rect 15210 2465 15216 2517
rect 15268 2465 15274 2517
rect 15210 2453 15274 2465
rect 15210 2401 15216 2453
rect 15268 2401 15274 2453
rect 15210 2394 15274 2401
rect 13269 2167 13315 2394
rect 13659 2167 13705 2394
rect 14049 2167 14095 2394
rect 14439 2167 14485 2394
rect 14829 2167 14875 2394
rect 15219 2167 15265 2394
rect 12891 2109 12897 2161
rect 12949 2109 12955 2161
rect 12891 2103 12955 2109
rect 13260 2161 13324 2167
rect 13260 2109 13266 2161
rect 13318 2109 13324 2161
rect 13260 2103 13324 2109
rect 13650 2161 13714 2167
rect 13650 2109 13656 2161
rect 13708 2109 13714 2161
rect 13650 2103 13714 2109
rect 14040 2161 14104 2167
rect 14040 2109 14046 2161
rect 14098 2109 14104 2161
rect 14040 2103 14104 2109
rect 14430 2161 14494 2167
rect 14430 2109 14436 2161
rect 14488 2109 14494 2161
rect 14430 2103 14494 2109
rect 14820 2161 14884 2167
rect 14820 2109 14826 2161
rect 14878 2109 14884 2161
rect 14820 2103 14884 2109
rect 15210 2161 15274 2167
rect 15210 2109 15216 2161
rect 15268 2109 15274 2161
rect 15210 2103 15274 2109
rect 15665 2161 15729 4065
rect 15665 2109 15671 2161
rect 15723 2109 15729 2161
rect 15665 2103 15729 2109
rect 13269 1884 13315 2103
rect 13659 1884 13705 2103
rect 14049 1884 14095 2103
rect 14439 1884 14485 2103
rect 14829 1884 14875 2103
rect 15219 1884 15265 2103
rect 13260 1865 13324 1884
rect 13260 1813 13266 1865
rect 13318 1813 13324 1865
rect 13260 1801 13324 1813
rect 13260 1749 13266 1801
rect 13318 1749 13324 1801
rect 13260 1737 13324 1749
rect 13260 1685 13266 1737
rect 13318 1685 13324 1737
rect 13260 1673 13324 1685
rect 13260 1621 13266 1673
rect 13318 1621 13324 1673
rect 13260 1609 13324 1621
rect 13260 1557 13266 1609
rect 13318 1557 13324 1609
rect 13260 1538 13324 1557
rect 13650 1865 13714 1884
rect 13650 1813 13656 1865
rect 13708 1813 13714 1865
rect 13650 1801 13714 1813
rect 13650 1749 13656 1801
rect 13708 1749 13714 1801
rect 13650 1737 13714 1749
rect 13650 1685 13656 1737
rect 13708 1685 13714 1737
rect 13650 1673 13714 1685
rect 13650 1621 13656 1673
rect 13708 1621 13714 1673
rect 13650 1609 13714 1621
rect 13650 1557 13656 1609
rect 13708 1557 13714 1609
rect 13650 1538 13714 1557
rect 14040 1865 14104 1884
rect 14040 1813 14046 1865
rect 14098 1813 14104 1865
rect 14040 1801 14104 1813
rect 14040 1749 14046 1801
rect 14098 1749 14104 1801
rect 14040 1737 14104 1749
rect 14040 1685 14046 1737
rect 14098 1685 14104 1737
rect 14040 1673 14104 1685
rect 14040 1621 14046 1673
rect 14098 1621 14104 1673
rect 14040 1609 14104 1621
rect 14040 1557 14046 1609
rect 14098 1557 14104 1609
rect 14040 1538 14104 1557
rect 14430 1865 14494 1884
rect 14430 1813 14436 1865
rect 14488 1813 14494 1865
rect 14430 1801 14494 1813
rect 14430 1749 14436 1801
rect 14488 1749 14494 1801
rect 14430 1737 14494 1749
rect 14430 1685 14436 1737
rect 14488 1685 14494 1737
rect 14430 1673 14494 1685
rect 14430 1621 14436 1673
rect 14488 1621 14494 1673
rect 14430 1609 14494 1621
rect 14430 1557 14436 1609
rect 14488 1557 14494 1609
rect 14430 1538 14494 1557
rect 14820 1865 14884 1884
rect 14820 1813 14826 1865
rect 14878 1813 14884 1865
rect 14820 1801 14884 1813
rect 14820 1749 14826 1801
rect 14878 1749 14884 1801
rect 14820 1737 14884 1749
rect 14820 1685 14826 1737
rect 14878 1685 14884 1737
rect 14820 1673 14884 1685
rect 14820 1621 14826 1673
rect 14878 1621 14884 1673
rect 14820 1609 14884 1621
rect 14820 1557 14826 1609
rect 14878 1557 14884 1609
rect 14820 1538 14884 1557
rect 15210 1865 15274 1884
rect 15210 1813 15216 1865
rect 15268 1813 15274 1865
rect 15210 1801 15274 1813
rect 15210 1749 15216 1801
rect 15268 1749 15274 1801
rect 15210 1737 15274 1749
rect 15210 1685 15216 1737
rect 15268 1685 15274 1737
rect 15210 1673 15274 1685
rect 15210 1621 15216 1673
rect 15268 1621 15274 1673
rect 15210 1609 15274 1621
rect 15210 1557 15216 1609
rect 15268 1557 15274 1609
rect 15210 1538 15274 1557
rect 13125 1191 13199 1213
rect 13125 1135 13134 1191
rect 13190 1135 13199 1191
rect 13125 1113 13199 1135
rect 13255 1191 13329 1213
rect 13255 1135 13264 1191
rect 13320 1135 13329 1191
rect 13255 1113 13329 1135
rect 13515 1191 13589 1213
rect 13515 1135 13524 1191
rect 13580 1135 13589 1191
rect 13515 1113 13589 1135
rect 13645 1191 13719 1213
rect 13645 1135 13654 1191
rect 13710 1135 13719 1191
rect 13645 1113 13719 1135
rect 13905 1191 13979 1213
rect 13905 1135 13914 1191
rect 13970 1135 13979 1191
rect 13905 1113 13979 1135
rect 14035 1191 14109 1213
rect 14035 1135 14044 1191
rect 14100 1135 14109 1191
rect 14035 1113 14109 1135
rect 14295 1191 14369 1213
rect 14295 1135 14304 1191
rect 14360 1135 14369 1191
rect 14295 1113 14369 1135
rect 14425 1191 14499 1213
rect 14425 1135 14434 1191
rect 14490 1135 14499 1191
rect 14425 1113 14499 1135
rect 14685 1191 14759 1213
rect 14685 1135 14694 1191
rect 14750 1135 14759 1191
rect 14685 1113 14759 1135
rect 14815 1191 14889 1213
rect 14815 1135 14824 1191
rect 14880 1135 14889 1191
rect 14815 1113 14889 1135
rect 15075 1191 15149 1213
rect 15075 1135 15084 1191
rect 15140 1135 15149 1191
rect 15075 1113 15149 1135
rect 15205 1191 15279 1213
rect 15205 1135 15214 1191
rect 15270 1135 15279 1191
rect 15205 1113 15279 1135
rect 15465 1191 15539 1213
rect 15465 1135 15474 1191
rect 15530 1135 15539 1191
rect 15465 1113 15539 1135
rect 24095 923 24149 5303
rect 24592 5217 24656 5303
rect 24592 5165 24598 5217
rect 24650 5165 24656 5217
rect 24592 5153 24656 5165
rect 24592 5101 24598 5153
rect 24650 5101 24656 5153
rect 24592 5089 24656 5101
rect 24592 5037 24598 5089
rect 24650 5037 24656 5089
rect 24592 5025 24656 5037
rect 24592 4973 24598 5025
rect 24650 4973 24656 5025
rect 24717 5091 24791 5113
rect 24717 5035 24726 5091
rect 24782 5035 24791 5091
rect 24717 5013 24791 5035
rect 24977 5091 25051 5113
rect 24977 5035 24986 5091
rect 25042 5035 25051 5091
rect 24977 5013 25051 5035
rect 25107 5091 25181 5113
rect 25107 5035 25116 5091
rect 25172 5035 25181 5091
rect 25107 5013 25181 5035
rect 25367 5091 25441 5113
rect 25367 5035 25376 5091
rect 25432 5035 25441 5091
rect 25367 5013 25441 5035
rect 25497 5091 25571 5113
rect 25497 5035 25506 5091
rect 25562 5035 25571 5091
rect 25497 5013 25571 5035
rect 25757 5091 25831 5113
rect 25757 5035 25766 5091
rect 25822 5035 25831 5091
rect 25757 5013 25831 5035
rect 25887 5091 25961 5113
rect 25887 5035 25896 5091
rect 25952 5035 25961 5091
rect 25887 5013 25961 5035
rect 26147 5091 26221 5113
rect 26147 5035 26156 5091
rect 26212 5035 26221 5091
rect 26147 5013 26221 5035
rect 26277 5091 26351 5113
rect 26277 5035 26286 5091
rect 26342 5035 26351 5091
rect 26277 5013 26351 5035
rect 26537 5091 26611 5113
rect 26537 5035 26546 5091
rect 26602 5035 26611 5091
rect 26537 5013 26611 5035
rect 26667 5091 26741 5113
rect 26667 5035 26676 5091
rect 26732 5035 26741 5091
rect 26667 5013 26741 5035
rect 24592 4961 24656 4973
rect 24592 4909 24598 4961
rect 24650 4909 24656 4961
rect 24483 4117 24547 4123
rect 24483 4065 24489 4117
rect 24541 4065 24547 4117
rect 24182 3960 24246 3961
rect 24182 3908 24188 3960
rect 24240 3908 24246 3960
rect 24182 3907 24246 3908
rect 24187 3405 24241 3907
rect 24177 3400 24251 3405
rect 24177 3344 24186 3400
rect 24242 3344 24251 3400
rect 24177 3339 24251 3344
rect 24187 2319 24241 3339
rect 24269 3274 24343 3279
rect 24269 3218 24278 3274
rect 24334 3218 24343 3274
rect 24269 3213 24343 3218
rect 24279 3013 24333 3213
rect 24269 3008 24343 3013
rect 24269 2952 24278 3008
rect 24334 2952 24343 3008
rect 24269 2947 24343 2952
rect 24182 2318 24246 2319
rect 24182 2266 24188 2318
rect 24240 2266 24246 2318
rect 24182 2265 24246 2266
rect 24483 2161 24547 4065
rect 24592 3477 24656 4909
rect 26799 4926 26999 4931
rect 26799 4870 26831 4926
rect 26887 4924 26911 4926
rect 26967 4925 26999 4926
rect 26967 4924 27110 4925
rect 26887 4872 26909 4924
rect 26967 4872 26973 4924
rect 27025 4872 27037 4924
rect 27089 4872 27110 4924
rect 26887 4870 26911 4872
rect 26967 4871 27110 4872
rect 26967 4870 26999 4871
rect 26799 4865 26999 4870
rect 26790 4781 26796 4833
rect 26848 4781 26854 4833
rect 24982 4669 25046 4688
rect 24982 4617 24988 4669
rect 25040 4617 25046 4669
rect 24982 4605 25046 4617
rect 24982 4553 24988 4605
rect 25040 4553 25046 4605
rect 24982 4541 25046 4553
rect 24982 4489 24988 4541
rect 25040 4489 25046 4541
rect 24982 4477 25046 4489
rect 24982 4425 24988 4477
rect 25040 4425 25046 4477
rect 24982 4413 25046 4425
rect 24982 4361 24988 4413
rect 25040 4361 25046 4413
rect 24982 4342 25046 4361
rect 25372 4669 25436 4688
rect 25372 4617 25378 4669
rect 25430 4617 25436 4669
rect 25372 4605 25436 4617
rect 25372 4553 25378 4605
rect 25430 4553 25436 4605
rect 25372 4541 25436 4553
rect 25372 4489 25378 4541
rect 25430 4489 25436 4541
rect 25372 4477 25436 4489
rect 25372 4425 25378 4477
rect 25430 4425 25436 4477
rect 25372 4413 25436 4425
rect 25372 4361 25378 4413
rect 25430 4361 25436 4413
rect 25372 4342 25436 4361
rect 25762 4669 25826 4688
rect 25762 4617 25768 4669
rect 25820 4617 25826 4669
rect 25762 4605 25826 4617
rect 25762 4553 25768 4605
rect 25820 4553 25826 4605
rect 25762 4541 25826 4553
rect 25762 4489 25768 4541
rect 25820 4489 25826 4541
rect 25762 4477 25826 4489
rect 25762 4425 25768 4477
rect 25820 4425 25826 4477
rect 25762 4413 25826 4425
rect 25762 4361 25768 4413
rect 25820 4361 25826 4413
rect 25762 4342 25826 4361
rect 26152 4669 26216 4688
rect 26152 4617 26158 4669
rect 26210 4617 26216 4669
rect 26152 4605 26216 4617
rect 26152 4553 26158 4605
rect 26210 4553 26216 4605
rect 26152 4541 26216 4553
rect 26152 4489 26158 4541
rect 26210 4489 26216 4541
rect 26152 4477 26216 4489
rect 26152 4425 26158 4477
rect 26210 4425 26216 4477
rect 26152 4413 26216 4425
rect 26152 4361 26158 4413
rect 26210 4361 26216 4413
rect 26152 4342 26216 4361
rect 26542 4669 26606 4688
rect 26542 4617 26548 4669
rect 26600 4617 26606 4669
rect 26542 4605 26606 4617
rect 26542 4553 26548 4605
rect 26600 4553 26606 4605
rect 26542 4541 26606 4553
rect 26542 4489 26548 4541
rect 26600 4489 26606 4541
rect 26542 4477 26606 4489
rect 26542 4425 26548 4477
rect 26600 4425 26606 4477
rect 26542 4413 26606 4425
rect 26542 4361 26548 4413
rect 26600 4361 26606 4413
rect 26797 4397 26837 4781
rect 26890 4685 26930 4865
rect 27067 4685 27107 4871
rect 26876 4633 26882 4685
rect 26934 4633 26940 4685
rect 27056 4633 27062 4685
rect 27114 4633 27120 4685
rect 26542 4342 26606 4361
rect 26786 4345 26792 4397
rect 26844 4345 26850 4397
rect 26965 4391 27031 4392
rect 24991 4123 25037 4342
rect 25381 4123 25427 4342
rect 25771 4123 25817 4342
rect 26161 4123 26207 4342
rect 26551 4123 26597 4342
rect 24982 4117 25046 4123
rect 24982 4065 24988 4117
rect 25040 4065 25046 4117
rect 24982 4059 25046 4065
rect 25372 4117 25436 4123
rect 25372 4065 25378 4117
rect 25430 4065 25436 4117
rect 25372 4059 25436 4065
rect 25762 4117 25826 4123
rect 25762 4065 25768 4117
rect 25820 4065 25826 4117
rect 25762 4059 25826 4065
rect 26152 4117 26216 4123
rect 26152 4065 26158 4117
rect 26210 4065 26216 4117
rect 26152 4059 26216 4065
rect 26542 4117 26606 4123
rect 26542 4065 26548 4117
rect 26600 4065 26606 4117
rect 26542 4059 26606 4065
rect 24991 3832 25037 4059
rect 25381 3832 25427 4059
rect 25771 3832 25817 4059
rect 26161 3832 26207 4059
rect 26551 3832 26597 4059
rect 24982 3825 25046 3832
rect 24982 3773 24988 3825
rect 25040 3773 25046 3825
rect 24982 3761 25046 3773
rect 24982 3709 24988 3761
rect 25040 3709 25046 3761
rect 24982 3702 25046 3709
rect 25112 3825 25176 3832
rect 25112 3773 25118 3825
rect 25170 3773 25176 3825
rect 25112 3761 25176 3773
rect 25112 3709 25118 3761
rect 25170 3709 25176 3761
rect 25112 3702 25176 3709
rect 25372 3825 25436 3832
rect 25372 3773 25378 3825
rect 25430 3773 25436 3825
rect 25372 3761 25436 3773
rect 25372 3709 25378 3761
rect 25430 3709 25436 3761
rect 25372 3702 25436 3709
rect 25502 3825 25566 3832
rect 25502 3773 25508 3825
rect 25560 3773 25566 3825
rect 25502 3761 25566 3773
rect 25502 3709 25508 3761
rect 25560 3709 25566 3761
rect 25502 3702 25566 3709
rect 25762 3825 25826 3832
rect 25762 3773 25768 3825
rect 25820 3773 25826 3825
rect 25762 3761 25826 3773
rect 25762 3709 25768 3761
rect 25820 3709 25826 3761
rect 25762 3702 25826 3709
rect 25892 3825 25956 3832
rect 25892 3773 25898 3825
rect 25950 3773 25956 3825
rect 25892 3761 25956 3773
rect 25892 3709 25898 3761
rect 25950 3709 25956 3761
rect 25892 3702 25956 3709
rect 26152 3825 26216 3832
rect 26152 3773 26158 3825
rect 26210 3773 26216 3825
rect 26152 3761 26216 3773
rect 26152 3709 26158 3761
rect 26210 3709 26216 3761
rect 26152 3702 26216 3709
rect 26282 3825 26346 3832
rect 26282 3773 26288 3825
rect 26340 3773 26346 3825
rect 26282 3761 26346 3773
rect 26282 3709 26288 3761
rect 26340 3709 26346 3761
rect 26282 3702 26346 3709
rect 26542 3825 26606 3832
rect 26542 3773 26548 3825
rect 26600 3773 26606 3825
rect 26542 3761 26606 3773
rect 26542 3709 26548 3761
rect 26600 3709 26606 3761
rect 26542 3702 26606 3709
rect 26672 3825 26736 3832
rect 26797 3829 26837 4345
rect 26965 4339 26972 4391
rect 27024 4339 27031 4391
rect 26965 4338 27031 4339
rect 27145 4391 27211 4392
rect 27145 4339 27152 4391
rect 27204 4339 27211 4391
rect 27145 4338 27211 4339
rect 26978 4296 27018 4338
rect 27158 4296 27198 4338
rect 27389 4297 27549 4302
rect 26965 4295 27031 4296
rect 26965 4243 26972 4295
rect 27024 4243 27031 4295
rect 26965 4242 27031 4243
rect 27145 4295 27211 4296
rect 27145 4243 27152 4295
rect 27204 4243 27211 4295
rect 27145 4242 27211 4243
rect 26978 3829 27018 4242
rect 27158 3829 27198 4242
rect 27389 4241 27401 4297
rect 27457 4295 27481 4297
rect 27463 4243 27475 4295
rect 27457 4241 27481 4243
rect 27537 4241 27549 4297
rect 27389 4236 27549 4241
rect 27257 4117 27321 4123
rect 27257 4065 27263 4117
rect 27315 4065 27321 4117
rect 26672 3773 26678 3825
rect 26730 3773 26736 3825
rect 26786 3777 26792 3829
rect 26844 3777 26850 3829
rect 26966 3777 26972 3829
rect 27024 3777 27030 3829
rect 27146 3777 27152 3829
rect 27204 3777 27210 3829
rect 26672 3761 26736 3773
rect 26672 3709 26678 3761
rect 26730 3709 26736 3761
rect 26672 3702 26736 3709
rect 26876 3705 26882 3757
rect 26934 3705 26940 3757
rect 27056 3705 27062 3757
rect 27114 3705 27120 3757
rect 24592 3425 24598 3477
rect 24650 3425 24656 3477
rect 25127 3469 25161 3702
rect 25517 3469 25551 3702
rect 25907 3469 25941 3702
rect 26297 3469 26331 3702
rect 26687 3469 26721 3702
rect 26886 3589 26926 3705
rect 27069 3595 27109 3705
rect 27059 3590 27229 3595
rect 27059 3589 27076 3590
rect 26886 3588 27076 3589
rect 26886 3536 26908 3588
rect 26960 3536 26972 3588
rect 27024 3536 27036 3588
rect 26886 3535 27076 3536
rect 26886 3533 26926 3535
rect 27059 3534 27076 3535
rect 27132 3534 27156 3590
rect 27212 3534 27229 3590
rect 27059 3529 27229 3534
rect 24592 3413 24656 3425
rect 24592 3361 24598 3413
rect 24650 3361 24656 3413
rect 24717 3447 24791 3469
rect 24717 3391 24726 3447
rect 24782 3391 24791 3447
rect 24717 3369 24791 3391
rect 24977 3447 25051 3469
rect 24977 3391 24986 3447
rect 25042 3391 25051 3447
rect 24977 3369 25051 3391
rect 25107 3447 25181 3469
rect 25107 3391 25116 3447
rect 25172 3391 25181 3447
rect 25107 3369 25181 3391
rect 25367 3447 25441 3469
rect 25367 3391 25376 3447
rect 25432 3391 25441 3447
rect 25367 3369 25441 3391
rect 25497 3447 25571 3469
rect 25497 3391 25506 3447
rect 25562 3391 25571 3447
rect 25497 3369 25571 3391
rect 25757 3447 25831 3469
rect 25757 3391 25766 3447
rect 25822 3391 25831 3447
rect 25757 3369 25831 3391
rect 25887 3447 25961 3469
rect 25887 3391 25896 3447
rect 25952 3391 25961 3447
rect 25887 3369 25961 3391
rect 26147 3447 26221 3469
rect 26147 3391 26156 3447
rect 26212 3391 26221 3447
rect 26147 3369 26221 3391
rect 26277 3447 26351 3469
rect 26277 3391 26286 3447
rect 26342 3391 26351 3447
rect 26277 3369 26351 3391
rect 26537 3447 26611 3469
rect 26537 3391 26546 3447
rect 26602 3391 26611 3447
rect 26537 3369 26611 3391
rect 26667 3447 26741 3469
rect 26667 3391 26676 3447
rect 26732 3391 26741 3447
rect 26667 3369 26741 3391
rect 24592 3354 24656 3361
rect 24584 3274 24658 3279
rect 24584 3218 24593 3274
rect 24649 3218 24658 3274
rect 24584 3213 24658 3218
rect 24912 3274 24986 3279
rect 24912 3218 24921 3274
rect 24977 3218 24986 3274
rect 24912 3213 24986 3218
rect 25302 3274 25376 3279
rect 25302 3218 25311 3274
rect 25367 3218 25376 3274
rect 25302 3213 25376 3218
rect 25692 3274 25766 3279
rect 25692 3218 25701 3274
rect 25757 3218 25766 3274
rect 25692 3213 25766 3218
rect 26082 3274 26156 3279
rect 26082 3218 26091 3274
rect 26147 3218 26156 3274
rect 26082 3213 26156 3218
rect 26472 3274 26546 3279
rect 26472 3218 26481 3274
rect 26537 3218 26546 3274
rect 26472 3213 26546 3218
rect 24849 3141 25049 3153
rect 24849 3139 24881 3141
rect 24937 3139 24961 3141
rect 25017 3139 25049 3141
rect 24849 3087 24859 3139
rect 25039 3087 25049 3139
rect 24849 3085 24881 3087
rect 24937 3085 24961 3087
rect 25017 3085 25049 3087
rect 24849 3073 25049 3085
rect 25629 3141 25829 3153
rect 25629 3139 25661 3141
rect 25717 3139 25741 3141
rect 25797 3139 25829 3141
rect 25629 3087 25639 3139
rect 25819 3087 25829 3139
rect 25629 3085 25661 3087
rect 25717 3085 25741 3087
rect 25797 3085 25829 3087
rect 25629 3073 25829 3085
rect 26409 3141 26609 3153
rect 26409 3139 26441 3141
rect 26497 3139 26521 3141
rect 26577 3139 26609 3141
rect 26409 3087 26419 3139
rect 26599 3087 26609 3139
rect 26409 3085 26441 3087
rect 26497 3085 26521 3087
rect 26577 3085 26609 3087
rect 26409 3073 26609 3085
rect 24912 3008 24986 3013
rect 24912 2952 24921 3008
rect 24977 2952 24986 3008
rect 24912 2947 24986 2952
rect 25302 3008 25376 3013
rect 25302 2952 25311 3008
rect 25367 2952 25376 3008
rect 25302 2947 25376 2952
rect 25692 3008 25766 3013
rect 25692 2952 25701 3008
rect 25757 2952 25766 3008
rect 25692 2947 25766 2952
rect 26082 3008 26156 3013
rect 26082 2952 26091 3008
rect 26147 2952 26156 3008
rect 26082 2947 26156 2952
rect 26472 3008 26546 3013
rect 26472 2952 26481 3008
rect 26537 2952 26546 3008
rect 26472 2947 26546 2952
rect 26862 3008 26936 3013
rect 26862 2952 26871 3008
rect 26927 2952 26936 3008
rect 26862 2947 26936 2952
rect 24717 2835 24791 2857
rect 24717 2779 24726 2835
rect 24782 2779 24791 2835
rect 24717 2757 24791 2779
rect 24847 2835 24921 2857
rect 24847 2779 24856 2835
rect 24912 2779 24921 2835
rect 24847 2757 24921 2779
rect 25107 2835 25181 2857
rect 25107 2779 25116 2835
rect 25172 2779 25181 2835
rect 25107 2757 25181 2779
rect 25237 2835 25311 2857
rect 25237 2779 25246 2835
rect 25302 2779 25311 2835
rect 25237 2757 25311 2779
rect 25497 2835 25571 2857
rect 25497 2779 25506 2835
rect 25562 2779 25571 2835
rect 25497 2757 25571 2779
rect 25627 2835 25701 2857
rect 25627 2779 25636 2835
rect 25692 2779 25701 2835
rect 25627 2757 25701 2779
rect 25887 2835 25961 2857
rect 25887 2779 25896 2835
rect 25952 2779 25961 2835
rect 25887 2757 25961 2779
rect 26017 2835 26091 2857
rect 26017 2779 26026 2835
rect 26082 2779 26091 2835
rect 26017 2757 26091 2779
rect 26277 2835 26351 2857
rect 26277 2779 26286 2835
rect 26342 2779 26351 2835
rect 26277 2757 26351 2779
rect 26407 2835 26481 2857
rect 26407 2779 26416 2835
rect 26472 2779 26481 2835
rect 26407 2757 26481 2779
rect 26667 2835 26741 2857
rect 26667 2779 26676 2835
rect 26732 2779 26741 2835
rect 26667 2757 26741 2779
rect 26797 2835 26871 2857
rect 26797 2779 26806 2835
rect 26862 2779 26871 2835
rect 26797 2757 26871 2779
rect 27057 2835 27131 2857
rect 27057 2779 27066 2835
rect 27122 2779 27131 2835
rect 27057 2757 27131 2779
rect 24737 2524 24771 2757
rect 25127 2524 25161 2757
rect 25517 2524 25551 2757
rect 25907 2524 25941 2757
rect 26297 2524 26331 2757
rect 26687 2524 26721 2757
rect 24722 2517 24786 2524
rect 24722 2465 24728 2517
rect 24780 2465 24786 2517
rect 24722 2453 24786 2465
rect 24722 2401 24728 2453
rect 24780 2401 24786 2453
rect 24722 2394 24786 2401
rect 24852 2517 24916 2524
rect 24852 2465 24858 2517
rect 24910 2465 24916 2517
rect 24852 2453 24916 2465
rect 24852 2401 24858 2453
rect 24910 2401 24916 2453
rect 24852 2394 24916 2401
rect 25112 2517 25176 2524
rect 25112 2465 25118 2517
rect 25170 2465 25176 2517
rect 25112 2453 25176 2465
rect 25112 2401 25118 2453
rect 25170 2401 25176 2453
rect 25112 2394 25176 2401
rect 25242 2517 25306 2524
rect 25242 2465 25248 2517
rect 25300 2465 25306 2517
rect 25242 2453 25306 2465
rect 25242 2401 25248 2453
rect 25300 2401 25306 2453
rect 25242 2394 25306 2401
rect 25502 2517 25566 2524
rect 25502 2465 25508 2517
rect 25560 2465 25566 2517
rect 25502 2453 25566 2465
rect 25502 2401 25508 2453
rect 25560 2401 25566 2453
rect 25502 2394 25566 2401
rect 25632 2517 25696 2524
rect 25632 2465 25638 2517
rect 25690 2465 25696 2517
rect 25632 2453 25696 2465
rect 25632 2401 25638 2453
rect 25690 2401 25696 2453
rect 25632 2394 25696 2401
rect 25892 2517 25956 2524
rect 25892 2465 25898 2517
rect 25950 2465 25956 2517
rect 25892 2453 25956 2465
rect 25892 2401 25898 2453
rect 25950 2401 25956 2453
rect 25892 2394 25956 2401
rect 26022 2517 26086 2524
rect 26022 2465 26028 2517
rect 26080 2465 26086 2517
rect 26022 2453 26086 2465
rect 26022 2401 26028 2453
rect 26080 2401 26086 2453
rect 26022 2394 26086 2401
rect 26282 2517 26346 2524
rect 26282 2465 26288 2517
rect 26340 2465 26346 2517
rect 26282 2453 26346 2465
rect 26282 2401 26288 2453
rect 26340 2401 26346 2453
rect 26282 2394 26346 2401
rect 26412 2517 26476 2524
rect 26412 2465 26418 2517
rect 26470 2465 26476 2517
rect 26412 2453 26476 2465
rect 26412 2401 26418 2453
rect 26470 2401 26476 2453
rect 26412 2394 26476 2401
rect 26672 2517 26736 2524
rect 26672 2465 26678 2517
rect 26730 2465 26736 2517
rect 26672 2453 26736 2465
rect 26672 2401 26678 2453
rect 26730 2401 26736 2453
rect 26672 2394 26736 2401
rect 26802 2517 26866 2524
rect 26802 2465 26808 2517
rect 26860 2465 26866 2517
rect 26802 2453 26866 2465
rect 26802 2401 26808 2453
rect 26860 2401 26866 2453
rect 26802 2394 26866 2401
rect 24861 2167 24907 2394
rect 25251 2167 25297 2394
rect 25641 2167 25687 2394
rect 26031 2167 26077 2394
rect 26421 2167 26467 2394
rect 26811 2167 26857 2394
rect 24483 2109 24489 2161
rect 24541 2109 24547 2161
rect 24483 2103 24547 2109
rect 24852 2161 24916 2167
rect 24852 2109 24858 2161
rect 24910 2109 24916 2161
rect 24852 2103 24916 2109
rect 25242 2161 25306 2167
rect 25242 2109 25248 2161
rect 25300 2109 25306 2161
rect 25242 2103 25306 2109
rect 25632 2161 25696 2167
rect 25632 2109 25638 2161
rect 25690 2109 25696 2161
rect 25632 2103 25696 2109
rect 26022 2161 26086 2167
rect 26022 2109 26028 2161
rect 26080 2109 26086 2161
rect 26022 2103 26086 2109
rect 26412 2161 26476 2167
rect 26412 2109 26418 2161
rect 26470 2109 26476 2161
rect 26412 2103 26476 2109
rect 26802 2161 26866 2167
rect 26802 2109 26808 2161
rect 26860 2109 26866 2161
rect 26802 2103 26866 2109
rect 27257 2161 27321 4065
rect 27257 2109 27263 2161
rect 27315 2109 27321 2161
rect 27257 2103 27321 2109
rect 24861 1884 24907 2103
rect 25251 1884 25297 2103
rect 25641 1884 25687 2103
rect 26031 1884 26077 2103
rect 26421 1884 26467 2103
rect 26811 1884 26857 2103
rect 24852 1865 24916 1884
rect 24852 1813 24858 1865
rect 24910 1813 24916 1865
rect 24852 1801 24916 1813
rect 24852 1749 24858 1801
rect 24910 1749 24916 1801
rect 24852 1737 24916 1749
rect 24852 1685 24858 1737
rect 24910 1685 24916 1737
rect 24852 1673 24916 1685
rect 24852 1621 24858 1673
rect 24910 1621 24916 1673
rect 24852 1609 24916 1621
rect 24852 1557 24858 1609
rect 24910 1557 24916 1609
rect 24852 1538 24916 1557
rect 25242 1865 25306 1884
rect 25242 1813 25248 1865
rect 25300 1813 25306 1865
rect 25242 1801 25306 1813
rect 25242 1749 25248 1801
rect 25300 1749 25306 1801
rect 25242 1737 25306 1749
rect 25242 1685 25248 1737
rect 25300 1685 25306 1737
rect 25242 1673 25306 1685
rect 25242 1621 25248 1673
rect 25300 1621 25306 1673
rect 25242 1609 25306 1621
rect 25242 1557 25248 1609
rect 25300 1557 25306 1609
rect 25242 1538 25306 1557
rect 25632 1865 25696 1884
rect 25632 1813 25638 1865
rect 25690 1813 25696 1865
rect 25632 1801 25696 1813
rect 25632 1749 25638 1801
rect 25690 1749 25696 1801
rect 25632 1737 25696 1749
rect 25632 1685 25638 1737
rect 25690 1685 25696 1737
rect 25632 1673 25696 1685
rect 25632 1621 25638 1673
rect 25690 1621 25696 1673
rect 25632 1609 25696 1621
rect 25632 1557 25638 1609
rect 25690 1557 25696 1609
rect 25632 1538 25696 1557
rect 26022 1865 26086 1884
rect 26022 1813 26028 1865
rect 26080 1813 26086 1865
rect 26022 1801 26086 1813
rect 26022 1749 26028 1801
rect 26080 1749 26086 1801
rect 26022 1737 26086 1749
rect 26022 1685 26028 1737
rect 26080 1685 26086 1737
rect 26022 1673 26086 1685
rect 26022 1621 26028 1673
rect 26080 1621 26086 1673
rect 26022 1609 26086 1621
rect 26022 1557 26028 1609
rect 26080 1557 26086 1609
rect 26022 1538 26086 1557
rect 26412 1865 26476 1884
rect 26412 1813 26418 1865
rect 26470 1813 26476 1865
rect 26412 1801 26476 1813
rect 26412 1749 26418 1801
rect 26470 1749 26476 1801
rect 26412 1737 26476 1749
rect 26412 1685 26418 1737
rect 26470 1685 26476 1737
rect 26412 1673 26476 1685
rect 26412 1621 26418 1673
rect 26470 1621 26476 1673
rect 26412 1609 26476 1621
rect 26412 1557 26418 1609
rect 26470 1557 26476 1609
rect 26412 1538 26476 1557
rect 26802 1865 26866 1884
rect 26802 1813 26808 1865
rect 26860 1813 26866 1865
rect 26802 1801 26866 1813
rect 26802 1749 26808 1801
rect 26860 1749 26866 1801
rect 26802 1737 26866 1749
rect 26802 1685 26808 1737
rect 26860 1685 26866 1737
rect 26802 1673 26866 1685
rect 26802 1621 26808 1673
rect 26860 1621 26866 1673
rect 26802 1609 26866 1621
rect 26802 1557 26808 1609
rect 26860 1557 26866 1609
rect 26802 1538 26866 1557
rect 24717 1191 24791 1213
rect 24717 1135 24726 1191
rect 24782 1135 24791 1191
rect 24717 1113 24791 1135
rect 24847 1191 24921 1213
rect 24847 1135 24856 1191
rect 24912 1135 24921 1191
rect 24847 1113 24921 1135
rect 25107 1191 25181 1213
rect 25107 1135 25116 1191
rect 25172 1135 25181 1191
rect 25107 1113 25181 1135
rect 25237 1191 25311 1213
rect 25237 1135 25246 1191
rect 25302 1135 25311 1191
rect 25237 1113 25311 1135
rect 25497 1191 25571 1213
rect 25497 1135 25506 1191
rect 25562 1135 25571 1191
rect 25497 1113 25571 1135
rect 25627 1191 25701 1213
rect 25627 1135 25636 1191
rect 25692 1135 25701 1191
rect 25627 1113 25701 1135
rect 25887 1191 25961 1213
rect 25887 1135 25896 1191
rect 25952 1135 25961 1191
rect 25887 1113 25961 1135
rect 26017 1191 26091 1213
rect 26017 1135 26026 1191
rect 26082 1135 26091 1191
rect 26017 1113 26091 1135
rect 26277 1191 26351 1213
rect 26277 1135 26286 1191
rect 26342 1135 26351 1191
rect 26277 1113 26351 1135
rect 26407 1191 26481 1213
rect 26407 1135 26416 1191
rect 26472 1135 26481 1191
rect 26407 1113 26481 1135
rect 26667 1191 26741 1213
rect 26667 1135 26676 1191
rect 26732 1135 26741 1191
rect 26667 1113 26741 1135
rect 26797 1191 26871 1213
rect 26797 1135 26806 1191
rect 26862 1135 26871 1191
rect 26797 1113 26871 1135
rect 27057 1191 27131 1213
rect 27057 1135 27066 1191
rect 27122 1135 27131 1191
rect 27057 1113 27131 1135
rect 12493 918 12567 923
rect 12493 862 12502 918
rect 12558 862 12567 918
rect 12493 857 12567 862
rect 13320 918 13394 923
rect 13320 862 13329 918
rect 13385 862 13394 918
rect 13320 857 13394 862
rect 13710 918 13784 923
rect 13710 862 13719 918
rect 13775 862 13784 918
rect 13710 857 13784 862
rect 14100 918 14174 923
rect 14100 862 14109 918
rect 14165 862 14174 918
rect 14100 857 14174 862
rect 14490 918 14564 923
rect 14490 862 14499 918
rect 14555 862 14564 918
rect 14490 857 14564 862
rect 14880 918 14954 923
rect 14880 862 14889 918
rect 14945 862 14954 918
rect 14880 857 14954 862
rect 15270 918 15344 923
rect 15270 862 15279 918
rect 15335 862 15344 918
rect 15270 857 15344 862
rect 24085 918 24159 923
rect 24085 862 24094 918
rect 24150 862 24159 918
rect 24085 857 24159 862
rect 24912 918 24986 923
rect 24912 862 24921 918
rect 24977 862 24986 918
rect 24912 857 24986 862
rect 25302 918 25376 923
rect 25302 862 25311 918
rect 25367 862 25376 918
rect 25302 857 25376 862
rect 25692 918 25766 923
rect 25692 862 25701 918
rect 25757 862 25766 918
rect 25692 857 25766 862
rect 26082 918 26156 923
rect 26082 862 26091 918
rect 26147 862 26156 918
rect 26082 857 26156 862
rect 26472 918 26546 923
rect 26472 862 26481 918
rect 26537 862 26546 918
rect 26472 857 26546 862
rect 26862 918 26936 923
rect 26862 862 26871 918
rect 26927 862 26936 918
rect 26862 857 26936 862
rect 12823 785 13023 797
rect 12823 783 12855 785
rect 12911 783 12935 785
rect 12991 783 13023 785
rect 12823 731 12833 783
rect 13013 731 13023 783
rect 12823 729 12855 731
rect 12911 729 12935 731
rect 12991 729 13023 731
rect 12823 717 13023 729
rect 13647 785 13847 797
rect 13647 783 13679 785
rect 13735 783 13759 785
rect 13815 783 13847 785
rect 13647 731 13657 783
rect 13837 731 13847 783
rect 13647 729 13679 731
rect 13735 729 13759 731
rect 13815 729 13847 731
rect 13647 717 13847 729
rect 14427 785 14627 797
rect 14427 783 14459 785
rect 14515 783 14539 785
rect 14595 783 14627 785
rect 14427 731 14437 783
rect 14617 731 14627 783
rect 14427 729 14459 731
rect 14515 729 14539 731
rect 14595 729 14627 731
rect 14427 717 14627 729
rect 15207 785 15407 797
rect 15207 783 15239 785
rect 15295 783 15319 785
rect 15375 783 15407 785
rect 15207 731 15217 783
rect 15397 731 15407 783
rect 15207 729 15239 731
rect 15295 729 15319 731
rect 15375 729 15407 731
rect 15207 717 15407 729
rect 24415 785 24615 797
rect 24415 783 24447 785
rect 24503 783 24527 785
rect 24583 783 24615 785
rect 24415 731 24425 783
rect 24605 731 24615 783
rect 24415 729 24447 731
rect 24503 729 24527 731
rect 24583 729 24615 731
rect 24415 717 24615 729
rect 25239 785 25439 797
rect 25239 783 25271 785
rect 25327 783 25351 785
rect 25407 783 25439 785
rect 25239 731 25249 783
rect 25429 731 25439 783
rect 25239 729 25271 731
rect 25327 729 25351 731
rect 25407 729 25439 731
rect 25239 717 25439 729
rect 26019 785 26219 797
rect 26019 783 26051 785
rect 26107 783 26131 785
rect 26187 783 26219 785
rect 26019 731 26029 783
rect 26209 731 26219 783
rect 26019 729 26051 731
rect 26107 729 26131 731
rect 26187 729 26219 731
rect 26019 717 26219 729
rect 26799 785 26999 797
rect 26799 783 26831 785
rect 26887 783 26911 785
rect 26967 783 26999 785
rect 26799 731 26809 783
rect 26989 731 26999 783
rect 26799 729 26831 731
rect 26887 729 26911 731
rect 26967 729 26999 731
rect 26799 717 26999 729
<< via2 >>
rect 12855 5495 12911 5497
rect 12935 5495 12991 5497
rect 12855 5443 12885 5495
rect 12885 5443 12897 5495
rect 12897 5443 12911 5495
rect 12935 5443 12949 5495
rect 12949 5443 12961 5495
rect 12961 5443 12991 5495
rect 12855 5441 12911 5443
rect 12935 5441 12991 5443
rect 13679 5495 13735 5497
rect 13759 5495 13815 5497
rect 13679 5443 13709 5495
rect 13709 5443 13721 5495
rect 13721 5443 13735 5495
rect 13759 5443 13773 5495
rect 13773 5443 13785 5495
rect 13785 5443 13815 5495
rect 13679 5441 13735 5443
rect 13759 5441 13815 5443
rect 14459 5495 14515 5497
rect 14539 5495 14595 5497
rect 14459 5443 14489 5495
rect 14489 5443 14501 5495
rect 14501 5443 14515 5495
rect 14539 5443 14553 5495
rect 14553 5443 14565 5495
rect 14565 5443 14595 5495
rect 14459 5441 14515 5443
rect 14539 5441 14595 5443
rect 15239 5495 15295 5497
rect 15319 5495 15375 5497
rect 15239 5443 15269 5495
rect 15269 5443 15281 5495
rect 15281 5443 15295 5495
rect 15319 5443 15333 5495
rect 15333 5443 15345 5495
rect 15345 5443 15375 5495
rect 15239 5441 15295 5443
rect 15319 5441 15375 5443
rect 24447 5495 24503 5497
rect 24527 5495 24583 5497
rect 24447 5443 24477 5495
rect 24477 5443 24489 5495
rect 24489 5443 24503 5495
rect 24527 5443 24541 5495
rect 24541 5443 24553 5495
rect 24553 5443 24583 5495
rect 24447 5441 24503 5443
rect 24527 5441 24583 5443
rect 25271 5495 25327 5497
rect 25351 5495 25407 5497
rect 25271 5443 25301 5495
rect 25301 5443 25313 5495
rect 25313 5443 25327 5495
rect 25351 5443 25365 5495
rect 25365 5443 25377 5495
rect 25377 5443 25407 5495
rect 25271 5441 25327 5443
rect 25351 5441 25407 5443
rect 26051 5495 26107 5497
rect 26131 5495 26187 5497
rect 26051 5443 26081 5495
rect 26081 5443 26093 5495
rect 26093 5443 26107 5495
rect 26131 5443 26145 5495
rect 26145 5443 26157 5495
rect 26157 5443 26187 5495
rect 26051 5441 26107 5443
rect 26131 5441 26187 5443
rect 26831 5495 26887 5497
rect 26911 5495 26967 5497
rect 26831 5443 26861 5495
rect 26861 5443 26873 5495
rect 26873 5443 26887 5495
rect 26911 5443 26925 5495
rect 26925 5443 26937 5495
rect 26937 5443 26967 5495
rect 26831 5441 26887 5443
rect 26911 5441 26967 5443
rect 12502 5362 12558 5364
rect 12502 5310 12504 5362
rect 12504 5310 12556 5362
rect 12556 5310 12558 5362
rect 12502 5308 12558 5310
rect 13039 5362 13095 5364
rect 13039 5310 13061 5362
rect 13061 5310 13073 5362
rect 13073 5310 13095 5362
rect 13039 5308 13095 5310
rect 13329 5362 13385 5364
rect 13329 5310 13331 5362
rect 13331 5310 13383 5362
rect 13383 5310 13385 5362
rect 13329 5308 13385 5310
rect 13719 5362 13775 5364
rect 13719 5310 13721 5362
rect 13721 5310 13773 5362
rect 13773 5310 13775 5362
rect 13719 5308 13775 5310
rect 14109 5362 14165 5364
rect 14109 5310 14111 5362
rect 14111 5310 14163 5362
rect 14163 5310 14165 5362
rect 14109 5308 14165 5310
rect 14499 5362 14555 5364
rect 14499 5310 14501 5362
rect 14501 5310 14553 5362
rect 14553 5310 14555 5362
rect 14499 5308 14555 5310
rect 14889 5362 14945 5364
rect 14889 5310 14891 5362
rect 14891 5310 14943 5362
rect 14943 5310 14945 5362
rect 14889 5308 14945 5310
rect 24094 5362 24150 5364
rect 24094 5310 24096 5362
rect 24096 5310 24148 5362
rect 24148 5310 24150 5362
rect 24094 5308 24150 5310
rect 24631 5362 24687 5364
rect 24631 5310 24653 5362
rect 24653 5310 24665 5362
rect 24665 5310 24687 5362
rect 24631 5308 24687 5310
rect 24921 5362 24977 5364
rect 24921 5310 24923 5362
rect 24923 5310 24975 5362
rect 24975 5310 24977 5362
rect 24921 5308 24977 5310
rect 25311 5362 25367 5364
rect 25311 5310 25313 5362
rect 25313 5310 25365 5362
rect 25365 5310 25367 5362
rect 25311 5308 25367 5310
rect 25701 5362 25757 5364
rect 25701 5310 25703 5362
rect 25703 5310 25755 5362
rect 25755 5310 25757 5362
rect 25701 5308 25757 5310
rect 26091 5362 26147 5364
rect 26091 5310 26093 5362
rect 26093 5310 26145 5362
rect 26145 5310 26147 5362
rect 26091 5308 26147 5310
rect 26481 5362 26537 5364
rect 26481 5310 26483 5362
rect 26483 5310 26535 5362
rect 26535 5310 26537 5362
rect 26481 5308 26537 5310
rect 13134 5089 13190 5091
rect 13134 5037 13136 5089
rect 13136 5037 13188 5089
rect 13188 5037 13190 5089
rect 13134 5035 13190 5037
rect 13394 5089 13450 5091
rect 13394 5037 13396 5089
rect 13396 5037 13448 5089
rect 13448 5037 13450 5089
rect 13394 5035 13450 5037
rect 13524 5089 13580 5091
rect 13524 5037 13526 5089
rect 13526 5037 13578 5089
rect 13578 5037 13580 5089
rect 13524 5035 13580 5037
rect 13784 5089 13840 5091
rect 13784 5037 13786 5089
rect 13786 5037 13838 5089
rect 13838 5037 13840 5089
rect 13784 5035 13840 5037
rect 13914 5089 13970 5091
rect 13914 5037 13916 5089
rect 13916 5037 13968 5089
rect 13968 5037 13970 5089
rect 13914 5035 13970 5037
rect 14174 5089 14230 5091
rect 14174 5037 14176 5089
rect 14176 5037 14228 5089
rect 14228 5037 14230 5089
rect 14174 5035 14230 5037
rect 14304 5089 14360 5091
rect 14304 5037 14306 5089
rect 14306 5037 14358 5089
rect 14358 5037 14360 5089
rect 14304 5035 14360 5037
rect 14564 5089 14620 5091
rect 14564 5037 14566 5089
rect 14566 5037 14618 5089
rect 14618 5037 14620 5089
rect 14564 5035 14620 5037
rect 14694 5089 14750 5091
rect 14694 5037 14696 5089
rect 14696 5037 14748 5089
rect 14748 5037 14750 5089
rect 14694 5035 14750 5037
rect 14954 5089 15010 5091
rect 14954 5037 14956 5089
rect 14956 5037 15008 5089
rect 15008 5037 15010 5089
rect 14954 5035 15010 5037
rect 15084 5089 15140 5091
rect 15084 5037 15086 5089
rect 15086 5037 15138 5089
rect 15138 5037 15140 5089
rect 15084 5035 15140 5037
rect 12594 3398 12650 3400
rect 12594 3346 12596 3398
rect 12596 3346 12648 3398
rect 12648 3346 12650 3398
rect 12594 3344 12650 3346
rect 12686 3272 12742 3274
rect 12686 3220 12688 3272
rect 12688 3220 12740 3272
rect 12740 3220 12742 3272
rect 12686 3218 12742 3220
rect 12686 3006 12742 3008
rect 12686 2954 12688 3006
rect 12688 2954 12740 3006
rect 12740 2954 12742 3006
rect 12686 2952 12742 2954
rect 15239 4870 15295 4926
rect 15319 4924 15375 4926
rect 15319 4872 15369 4924
rect 15369 4872 15375 4924
rect 15319 4870 15375 4872
rect 15809 4295 15865 4297
rect 15889 4295 15945 4297
rect 15809 4243 15819 4295
rect 15819 4243 15865 4295
rect 15889 4243 15935 4295
rect 15935 4243 15945 4295
rect 15809 4241 15865 4243
rect 15889 4241 15945 4243
rect 15484 3588 15540 3590
rect 15484 3536 15496 3588
rect 15496 3536 15540 3588
rect 15484 3534 15540 3536
rect 15564 3534 15620 3590
rect 13134 3445 13190 3447
rect 13134 3393 13136 3445
rect 13136 3393 13188 3445
rect 13188 3393 13190 3445
rect 13134 3391 13190 3393
rect 13394 3445 13450 3447
rect 13394 3393 13396 3445
rect 13396 3393 13448 3445
rect 13448 3393 13450 3445
rect 13394 3391 13450 3393
rect 13524 3445 13580 3447
rect 13524 3393 13526 3445
rect 13526 3393 13578 3445
rect 13578 3393 13580 3445
rect 13524 3391 13580 3393
rect 13784 3445 13840 3447
rect 13784 3393 13786 3445
rect 13786 3393 13838 3445
rect 13838 3393 13840 3445
rect 13784 3391 13840 3393
rect 13914 3445 13970 3447
rect 13914 3393 13916 3445
rect 13916 3393 13968 3445
rect 13968 3393 13970 3445
rect 13914 3391 13970 3393
rect 14174 3445 14230 3447
rect 14174 3393 14176 3445
rect 14176 3393 14228 3445
rect 14228 3393 14230 3445
rect 14174 3391 14230 3393
rect 14304 3445 14360 3447
rect 14304 3393 14306 3445
rect 14306 3393 14358 3445
rect 14358 3393 14360 3445
rect 14304 3391 14360 3393
rect 14564 3445 14620 3447
rect 14564 3393 14566 3445
rect 14566 3393 14618 3445
rect 14618 3393 14620 3445
rect 14564 3391 14620 3393
rect 14694 3445 14750 3447
rect 14694 3393 14696 3445
rect 14696 3393 14748 3445
rect 14748 3393 14750 3445
rect 14694 3391 14750 3393
rect 14954 3445 15010 3447
rect 14954 3393 14956 3445
rect 14956 3393 15008 3445
rect 15008 3393 15010 3445
rect 14954 3391 15010 3393
rect 15084 3445 15140 3447
rect 15084 3393 15086 3445
rect 15086 3393 15138 3445
rect 15138 3393 15140 3445
rect 15084 3391 15140 3393
rect 13001 3272 13057 3274
rect 13001 3220 13003 3272
rect 13003 3220 13055 3272
rect 13055 3220 13057 3272
rect 13001 3218 13057 3220
rect 13329 3272 13385 3274
rect 13329 3220 13331 3272
rect 13331 3220 13383 3272
rect 13383 3220 13385 3272
rect 13329 3218 13385 3220
rect 13719 3272 13775 3274
rect 13719 3220 13721 3272
rect 13721 3220 13773 3272
rect 13773 3220 13775 3272
rect 13719 3218 13775 3220
rect 14109 3272 14165 3274
rect 14109 3220 14111 3272
rect 14111 3220 14163 3272
rect 14163 3220 14165 3272
rect 14109 3218 14165 3220
rect 14499 3272 14555 3274
rect 14499 3220 14501 3272
rect 14501 3220 14553 3272
rect 14553 3220 14555 3272
rect 14499 3218 14555 3220
rect 14889 3272 14945 3274
rect 14889 3220 14891 3272
rect 14891 3220 14943 3272
rect 14943 3220 14945 3272
rect 14889 3218 14945 3220
rect 13289 3139 13345 3141
rect 13369 3139 13425 3141
rect 13289 3087 13319 3139
rect 13319 3087 13331 3139
rect 13331 3087 13345 3139
rect 13369 3087 13383 3139
rect 13383 3087 13395 3139
rect 13395 3087 13425 3139
rect 13289 3085 13345 3087
rect 13369 3085 13425 3087
rect 14069 3139 14125 3141
rect 14149 3139 14205 3141
rect 14069 3087 14099 3139
rect 14099 3087 14111 3139
rect 14111 3087 14125 3139
rect 14149 3087 14163 3139
rect 14163 3087 14175 3139
rect 14175 3087 14205 3139
rect 14069 3085 14125 3087
rect 14149 3085 14205 3087
rect 14849 3139 14905 3141
rect 14929 3139 14985 3141
rect 14849 3087 14879 3139
rect 14879 3087 14891 3139
rect 14891 3087 14905 3139
rect 14929 3087 14943 3139
rect 14943 3087 14955 3139
rect 14955 3087 14985 3139
rect 14849 3085 14905 3087
rect 14929 3085 14985 3087
rect 13329 3006 13385 3008
rect 13329 2954 13331 3006
rect 13331 2954 13383 3006
rect 13383 2954 13385 3006
rect 13329 2952 13385 2954
rect 13719 3006 13775 3008
rect 13719 2954 13721 3006
rect 13721 2954 13773 3006
rect 13773 2954 13775 3006
rect 13719 2952 13775 2954
rect 14109 3006 14165 3008
rect 14109 2954 14111 3006
rect 14111 2954 14163 3006
rect 14163 2954 14165 3006
rect 14109 2952 14165 2954
rect 14499 3006 14555 3008
rect 14499 2954 14501 3006
rect 14501 2954 14553 3006
rect 14553 2954 14555 3006
rect 14499 2952 14555 2954
rect 14889 3006 14945 3008
rect 14889 2954 14891 3006
rect 14891 2954 14943 3006
rect 14943 2954 14945 3006
rect 14889 2952 14945 2954
rect 15279 3006 15335 3008
rect 15279 2954 15281 3006
rect 15281 2954 15333 3006
rect 15333 2954 15335 3006
rect 15279 2952 15335 2954
rect 13134 2833 13190 2835
rect 13134 2781 13136 2833
rect 13136 2781 13188 2833
rect 13188 2781 13190 2833
rect 13134 2779 13190 2781
rect 13264 2833 13320 2835
rect 13264 2781 13266 2833
rect 13266 2781 13318 2833
rect 13318 2781 13320 2833
rect 13264 2779 13320 2781
rect 13524 2833 13580 2835
rect 13524 2781 13526 2833
rect 13526 2781 13578 2833
rect 13578 2781 13580 2833
rect 13524 2779 13580 2781
rect 13654 2833 13710 2835
rect 13654 2781 13656 2833
rect 13656 2781 13708 2833
rect 13708 2781 13710 2833
rect 13654 2779 13710 2781
rect 13914 2833 13970 2835
rect 13914 2781 13916 2833
rect 13916 2781 13968 2833
rect 13968 2781 13970 2833
rect 13914 2779 13970 2781
rect 14044 2833 14100 2835
rect 14044 2781 14046 2833
rect 14046 2781 14098 2833
rect 14098 2781 14100 2833
rect 14044 2779 14100 2781
rect 14304 2833 14360 2835
rect 14304 2781 14306 2833
rect 14306 2781 14358 2833
rect 14358 2781 14360 2833
rect 14304 2779 14360 2781
rect 14434 2833 14490 2835
rect 14434 2781 14436 2833
rect 14436 2781 14488 2833
rect 14488 2781 14490 2833
rect 14434 2779 14490 2781
rect 14694 2833 14750 2835
rect 14694 2781 14696 2833
rect 14696 2781 14748 2833
rect 14748 2781 14750 2833
rect 14694 2779 14750 2781
rect 14824 2833 14880 2835
rect 14824 2781 14826 2833
rect 14826 2781 14878 2833
rect 14878 2781 14880 2833
rect 14824 2779 14880 2781
rect 15084 2833 15140 2835
rect 15084 2781 15086 2833
rect 15086 2781 15138 2833
rect 15138 2781 15140 2833
rect 15084 2779 15140 2781
rect 15214 2833 15270 2835
rect 15214 2781 15216 2833
rect 15216 2781 15268 2833
rect 15268 2781 15270 2833
rect 15214 2779 15270 2781
rect 15474 2833 15530 2835
rect 15474 2781 15476 2833
rect 15476 2781 15528 2833
rect 15528 2781 15530 2833
rect 15474 2779 15530 2781
rect 13134 1189 13190 1191
rect 13134 1137 13136 1189
rect 13136 1137 13188 1189
rect 13188 1137 13190 1189
rect 13134 1135 13190 1137
rect 13264 1189 13320 1191
rect 13264 1137 13266 1189
rect 13266 1137 13318 1189
rect 13318 1137 13320 1189
rect 13264 1135 13320 1137
rect 13524 1189 13580 1191
rect 13524 1137 13526 1189
rect 13526 1137 13578 1189
rect 13578 1137 13580 1189
rect 13524 1135 13580 1137
rect 13654 1189 13710 1191
rect 13654 1137 13656 1189
rect 13656 1137 13708 1189
rect 13708 1137 13710 1189
rect 13654 1135 13710 1137
rect 13914 1189 13970 1191
rect 13914 1137 13916 1189
rect 13916 1137 13968 1189
rect 13968 1137 13970 1189
rect 13914 1135 13970 1137
rect 14044 1189 14100 1191
rect 14044 1137 14046 1189
rect 14046 1137 14098 1189
rect 14098 1137 14100 1189
rect 14044 1135 14100 1137
rect 14304 1189 14360 1191
rect 14304 1137 14306 1189
rect 14306 1137 14358 1189
rect 14358 1137 14360 1189
rect 14304 1135 14360 1137
rect 14434 1189 14490 1191
rect 14434 1137 14436 1189
rect 14436 1137 14488 1189
rect 14488 1137 14490 1189
rect 14434 1135 14490 1137
rect 14694 1189 14750 1191
rect 14694 1137 14696 1189
rect 14696 1137 14748 1189
rect 14748 1137 14750 1189
rect 14694 1135 14750 1137
rect 14824 1189 14880 1191
rect 14824 1137 14826 1189
rect 14826 1137 14878 1189
rect 14878 1137 14880 1189
rect 14824 1135 14880 1137
rect 15084 1189 15140 1191
rect 15084 1137 15086 1189
rect 15086 1137 15138 1189
rect 15138 1137 15140 1189
rect 15084 1135 15140 1137
rect 15214 1189 15270 1191
rect 15214 1137 15216 1189
rect 15216 1137 15268 1189
rect 15268 1137 15270 1189
rect 15214 1135 15270 1137
rect 15474 1189 15530 1191
rect 15474 1137 15476 1189
rect 15476 1137 15528 1189
rect 15528 1137 15530 1189
rect 15474 1135 15530 1137
rect 24726 5089 24782 5091
rect 24726 5037 24728 5089
rect 24728 5037 24780 5089
rect 24780 5037 24782 5089
rect 24726 5035 24782 5037
rect 24986 5089 25042 5091
rect 24986 5037 24988 5089
rect 24988 5037 25040 5089
rect 25040 5037 25042 5089
rect 24986 5035 25042 5037
rect 25116 5089 25172 5091
rect 25116 5037 25118 5089
rect 25118 5037 25170 5089
rect 25170 5037 25172 5089
rect 25116 5035 25172 5037
rect 25376 5089 25432 5091
rect 25376 5037 25378 5089
rect 25378 5037 25430 5089
rect 25430 5037 25432 5089
rect 25376 5035 25432 5037
rect 25506 5089 25562 5091
rect 25506 5037 25508 5089
rect 25508 5037 25560 5089
rect 25560 5037 25562 5089
rect 25506 5035 25562 5037
rect 25766 5089 25822 5091
rect 25766 5037 25768 5089
rect 25768 5037 25820 5089
rect 25820 5037 25822 5089
rect 25766 5035 25822 5037
rect 25896 5089 25952 5091
rect 25896 5037 25898 5089
rect 25898 5037 25950 5089
rect 25950 5037 25952 5089
rect 25896 5035 25952 5037
rect 26156 5089 26212 5091
rect 26156 5037 26158 5089
rect 26158 5037 26210 5089
rect 26210 5037 26212 5089
rect 26156 5035 26212 5037
rect 26286 5089 26342 5091
rect 26286 5037 26288 5089
rect 26288 5037 26340 5089
rect 26340 5037 26342 5089
rect 26286 5035 26342 5037
rect 26546 5089 26602 5091
rect 26546 5037 26548 5089
rect 26548 5037 26600 5089
rect 26600 5037 26602 5089
rect 26546 5035 26602 5037
rect 26676 5089 26732 5091
rect 26676 5037 26678 5089
rect 26678 5037 26730 5089
rect 26730 5037 26732 5089
rect 26676 5035 26732 5037
rect 24186 3398 24242 3400
rect 24186 3346 24188 3398
rect 24188 3346 24240 3398
rect 24240 3346 24242 3398
rect 24186 3344 24242 3346
rect 24278 3272 24334 3274
rect 24278 3220 24280 3272
rect 24280 3220 24332 3272
rect 24332 3220 24334 3272
rect 24278 3218 24334 3220
rect 24278 3006 24334 3008
rect 24278 2954 24280 3006
rect 24280 2954 24332 3006
rect 24332 2954 24334 3006
rect 24278 2952 24334 2954
rect 26831 4870 26887 4926
rect 26911 4924 26967 4926
rect 26911 4872 26961 4924
rect 26961 4872 26967 4924
rect 26911 4870 26967 4872
rect 27401 4295 27457 4297
rect 27481 4295 27537 4297
rect 27401 4243 27411 4295
rect 27411 4243 27457 4295
rect 27481 4243 27527 4295
rect 27527 4243 27537 4295
rect 27401 4241 27457 4243
rect 27481 4241 27537 4243
rect 27076 3588 27132 3590
rect 27076 3536 27088 3588
rect 27088 3536 27132 3588
rect 27076 3534 27132 3536
rect 27156 3534 27212 3590
rect 24726 3445 24782 3447
rect 24726 3393 24728 3445
rect 24728 3393 24780 3445
rect 24780 3393 24782 3445
rect 24726 3391 24782 3393
rect 24986 3445 25042 3447
rect 24986 3393 24988 3445
rect 24988 3393 25040 3445
rect 25040 3393 25042 3445
rect 24986 3391 25042 3393
rect 25116 3445 25172 3447
rect 25116 3393 25118 3445
rect 25118 3393 25170 3445
rect 25170 3393 25172 3445
rect 25116 3391 25172 3393
rect 25376 3445 25432 3447
rect 25376 3393 25378 3445
rect 25378 3393 25430 3445
rect 25430 3393 25432 3445
rect 25376 3391 25432 3393
rect 25506 3445 25562 3447
rect 25506 3393 25508 3445
rect 25508 3393 25560 3445
rect 25560 3393 25562 3445
rect 25506 3391 25562 3393
rect 25766 3445 25822 3447
rect 25766 3393 25768 3445
rect 25768 3393 25820 3445
rect 25820 3393 25822 3445
rect 25766 3391 25822 3393
rect 25896 3445 25952 3447
rect 25896 3393 25898 3445
rect 25898 3393 25950 3445
rect 25950 3393 25952 3445
rect 25896 3391 25952 3393
rect 26156 3445 26212 3447
rect 26156 3393 26158 3445
rect 26158 3393 26210 3445
rect 26210 3393 26212 3445
rect 26156 3391 26212 3393
rect 26286 3445 26342 3447
rect 26286 3393 26288 3445
rect 26288 3393 26340 3445
rect 26340 3393 26342 3445
rect 26286 3391 26342 3393
rect 26546 3445 26602 3447
rect 26546 3393 26548 3445
rect 26548 3393 26600 3445
rect 26600 3393 26602 3445
rect 26546 3391 26602 3393
rect 26676 3445 26732 3447
rect 26676 3393 26678 3445
rect 26678 3393 26730 3445
rect 26730 3393 26732 3445
rect 26676 3391 26732 3393
rect 24593 3272 24649 3274
rect 24593 3220 24595 3272
rect 24595 3220 24647 3272
rect 24647 3220 24649 3272
rect 24593 3218 24649 3220
rect 24921 3272 24977 3274
rect 24921 3220 24923 3272
rect 24923 3220 24975 3272
rect 24975 3220 24977 3272
rect 24921 3218 24977 3220
rect 25311 3272 25367 3274
rect 25311 3220 25313 3272
rect 25313 3220 25365 3272
rect 25365 3220 25367 3272
rect 25311 3218 25367 3220
rect 25701 3272 25757 3274
rect 25701 3220 25703 3272
rect 25703 3220 25755 3272
rect 25755 3220 25757 3272
rect 25701 3218 25757 3220
rect 26091 3272 26147 3274
rect 26091 3220 26093 3272
rect 26093 3220 26145 3272
rect 26145 3220 26147 3272
rect 26091 3218 26147 3220
rect 26481 3272 26537 3274
rect 26481 3220 26483 3272
rect 26483 3220 26535 3272
rect 26535 3220 26537 3272
rect 26481 3218 26537 3220
rect 24881 3139 24937 3141
rect 24961 3139 25017 3141
rect 24881 3087 24911 3139
rect 24911 3087 24923 3139
rect 24923 3087 24937 3139
rect 24961 3087 24975 3139
rect 24975 3087 24987 3139
rect 24987 3087 25017 3139
rect 24881 3085 24937 3087
rect 24961 3085 25017 3087
rect 25661 3139 25717 3141
rect 25741 3139 25797 3141
rect 25661 3087 25691 3139
rect 25691 3087 25703 3139
rect 25703 3087 25717 3139
rect 25741 3087 25755 3139
rect 25755 3087 25767 3139
rect 25767 3087 25797 3139
rect 25661 3085 25717 3087
rect 25741 3085 25797 3087
rect 26441 3139 26497 3141
rect 26521 3139 26577 3141
rect 26441 3087 26471 3139
rect 26471 3087 26483 3139
rect 26483 3087 26497 3139
rect 26521 3087 26535 3139
rect 26535 3087 26547 3139
rect 26547 3087 26577 3139
rect 26441 3085 26497 3087
rect 26521 3085 26577 3087
rect 24921 3006 24977 3008
rect 24921 2954 24923 3006
rect 24923 2954 24975 3006
rect 24975 2954 24977 3006
rect 24921 2952 24977 2954
rect 25311 3006 25367 3008
rect 25311 2954 25313 3006
rect 25313 2954 25365 3006
rect 25365 2954 25367 3006
rect 25311 2952 25367 2954
rect 25701 3006 25757 3008
rect 25701 2954 25703 3006
rect 25703 2954 25755 3006
rect 25755 2954 25757 3006
rect 25701 2952 25757 2954
rect 26091 3006 26147 3008
rect 26091 2954 26093 3006
rect 26093 2954 26145 3006
rect 26145 2954 26147 3006
rect 26091 2952 26147 2954
rect 26481 3006 26537 3008
rect 26481 2954 26483 3006
rect 26483 2954 26535 3006
rect 26535 2954 26537 3006
rect 26481 2952 26537 2954
rect 26871 3006 26927 3008
rect 26871 2954 26873 3006
rect 26873 2954 26925 3006
rect 26925 2954 26927 3006
rect 26871 2952 26927 2954
rect 24726 2833 24782 2835
rect 24726 2781 24728 2833
rect 24728 2781 24780 2833
rect 24780 2781 24782 2833
rect 24726 2779 24782 2781
rect 24856 2833 24912 2835
rect 24856 2781 24858 2833
rect 24858 2781 24910 2833
rect 24910 2781 24912 2833
rect 24856 2779 24912 2781
rect 25116 2833 25172 2835
rect 25116 2781 25118 2833
rect 25118 2781 25170 2833
rect 25170 2781 25172 2833
rect 25116 2779 25172 2781
rect 25246 2833 25302 2835
rect 25246 2781 25248 2833
rect 25248 2781 25300 2833
rect 25300 2781 25302 2833
rect 25246 2779 25302 2781
rect 25506 2833 25562 2835
rect 25506 2781 25508 2833
rect 25508 2781 25560 2833
rect 25560 2781 25562 2833
rect 25506 2779 25562 2781
rect 25636 2833 25692 2835
rect 25636 2781 25638 2833
rect 25638 2781 25690 2833
rect 25690 2781 25692 2833
rect 25636 2779 25692 2781
rect 25896 2833 25952 2835
rect 25896 2781 25898 2833
rect 25898 2781 25950 2833
rect 25950 2781 25952 2833
rect 25896 2779 25952 2781
rect 26026 2833 26082 2835
rect 26026 2781 26028 2833
rect 26028 2781 26080 2833
rect 26080 2781 26082 2833
rect 26026 2779 26082 2781
rect 26286 2833 26342 2835
rect 26286 2781 26288 2833
rect 26288 2781 26340 2833
rect 26340 2781 26342 2833
rect 26286 2779 26342 2781
rect 26416 2833 26472 2835
rect 26416 2781 26418 2833
rect 26418 2781 26470 2833
rect 26470 2781 26472 2833
rect 26416 2779 26472 2781
rect 26676 2833 26732 2835
rect 26676 2781 26678 2833
rect 26678 2781 26730 2833
rect 26730 2781 26732 2833
rect 26676 2779 26732 2781
rect 26806 2833 26862 2835
rect 26806 2781 26808 2833
rect 26808 2781 26860 2833
rect 26860 2781 26862 2833
rect 26806 2779 26862 2781
rect 27066 2833 27122 2835
rect 27066 2781 27068 2833
rect 27068 2781 27120 2833
rect 27120 2781 27122 2833
rect 27066 2779 27122 2781
rect 24726 1189 24782 1191
rect 24726 1137 24728 1189
rect 24728 1137 24780 1189
rect 24780 1137 24782 1189
rect 24726 1135 24782 1137
rect 24856 1189 24912 1191
rect 24856 1137 24858 1189
rect 24858 1137 24910 1189
rect 24910 1137 24912 1189
rect 24856 1135 24912 1137
rect 25116 1189 25172 1191
rect 25116 1137 25118 1189
rect 25118 1137 25170 1189
rect 25170 1137 25172 1189
rect 25116 1135 25172 1137
rect 25246 1189 25302 1191
rect 25246 1137 25248 1189
rect 25248 1137 25300 1189
rect 25300 1137 25302 1189
rect 25246 1135 25302 1137
rect 25506 1189 25562 1191
rect 25506 1137 25508 1189
rect 25508 1137 25560 1189
rect 25560 1137 25562 1189
rect 25506 1135 25562 1137
rect 25636 1189 25692 1191
rect 25636 1137 25638 1189
rect 25638 1137 25690 1189
rect 25690 1137 25692 1189
rect 25636 1135 25692 1137
rect 25896 1189 25952 1191
rect 25896 1137 25898 1189
rect 25898 1137 25950 1189
rect 25950 1137 25952 1189
rect 25896 1135 25952 1137
rect 26026 1189 26082 1191
rect 26026 1137 26028 1189
rect 26028 1137 26080 1189
rect 26080 1137 26082 1189
rect 26026 1135 26082 1137
rect 26286 1189 26342 1191
rect 26286 1137 26288 1189
rect 26288 1137 26340 1189
rect 26340 1137 26342 1189
rect 26286 1135 26342 1137
rect 26416 1189 26472 1191
rect 26416 1137 26418 1189
rect 26418 1137 26470 1189
rect 26470 1137 26472 1189
rect 26416 1135 26472 1137
rect 26676 1189 26732 1191
rect 26676 1137 26678 1189
rect 26678 1137 26730 1189
rect 26730 1137 26732 1189
rect 26676 1135 26732 1137
rect 26806 1189 26862 1191
rect 26806 1137 26808 1189
rect 26808 1137 26860 1189
rect 26860 1137 26862 1189
rect 26806 1135 26862 1137
rect 27066 1189 27122 1191
rect 27066 1137 27068 1189
rect 27068 1137 27120 1189
rect 27120 1137 27122 1189
rect 27066 1135 27122 1137
rect 12502 916 12558 918
rect 12502 864 12504 916
rect 12504 864 12556 916
rect 12556 864 12558 916
rect 12502 862 12558 864
rect 13329 916 13385 918
rect 13329 864 13331 916
rect 13331 864 13383 916
rect 13383 864 13385 916
rect 13329 862 13385 864
rect 13719 916 13775 918
rect 13719 864 13721 916
rect 13721 864 13773 916
rect 13773 864 13775 916
rect 13719 862 13775 864
rect 14109 916 14165 918
rect 14109 864 14111 916
rect 14111 864 14163 916
rect 14163 864 14165 916
rect 14109 862 14165 864
rect 14499 916 14555 918
rect 14499 864 14501 916
rect 14501 864 14553 916
rect 14553 864 14555 916
rect 14499 862 14555 864
rect 14889 916 14945 918
rect 14889 864 14891 916
rect 14891 864 14943 916
rect 14943 864 14945 916
rect 14889 862 14945 864
rect 15279 916 15335 918
rect 15279 864 15281 916
rect 15281 864 15333 916
rect 15333 864 15335 916
rect 15279 862 15335 864
rect 24094 916 24150 918
rect 24094 864 24096 916
rect 24096 864 24148 916
rect 24148 864 24150 916
rect 24094 862 24150 864
rect 24921 916 24977 918
rect 24921 864 24923 916
rect 24923 864 24975 916
rect 24975 864 24977 916
rect 24921 862 24977 864
rect 25311 916 25367 918
rect 25311 864 25313 916
rect 25313 864 25365 916
rect 25365 864 25367 916
rect 25311 862 25367 864
rect 25701 916 25757 918
rect 25701 864 25703 916
rect 25703 864 25755 916
rect 25755 864 25757 916
rect 25701 862 25757 864
rect 26091 916 26147 918
rect 26091 864 26093 916
rect 26093 864 26145 916
rect 26145 864 26147 916
rect 26091 862 26147 864
rect 26481 916 26537 918
rect 26481 864 26483 916
rect 26483 864 26535 916
rect 26535 864 26537 916
rect 26481 862 26537 864
rect 26871 916 26927 918
rect 26871 864 26873 916
rect 26873 864 26925 916
rect 26925 864 26927 916
rect 26871 862 26927 864
rect 12855 783 12911 785
rect 12935 783 12991 785
rect 12855 731 12885 783
rect 12885 731 12897 783
rect 12897 731 12911 783
rect 12935 731 12949 783
rect 12949 731 12961 783
rect 12961 731 12991 783
rect 12855 729 12911 731
rect 12935 729 12991 731
rect 13679 783 13735 785
rect 13759 783 13815 785
rect 13679 731 13709 783
rect 13709 731 13721 783
rect 13721 731 13735 783
rect 13759 731 13773 783
rect 13773 731 13785 783
rect 13785 731 13815 783
rect 13679 729 13735 731
rect 13759 729 13815 731
rect 14459 783 14515 785
rect 14539 783 14595 785
rect 14459 731 14489 783
rect 14489 731 14501 783
rect 14501 731 14515 783
rect 14539 731 14553 783
rect 14553 731 14565 783
rect 14565 731 14595 783
rect 14459 729 14515 731
rect 14539 729 14595 731
rect 15239 783 15295 785
rect 15319 783 15375 785
rect 15239 731 15269 783
rect 15269 731 15281 783
rect 15281 731 15295 783
rect 15319 731 15333 783
rect 15333 731 15345 783
rect 15345 731 15375 783
rect 15239 729 15295 731
rect 15319 729 15375 731
rect 24447 783 24503 785
rect 24527 783 24583 785
rect 24447 731 24477 783
rect 24477 731 24489 783
rect 24489 731 24503 783
rect 24527 731 24541 783
rect 24541 731 24553 783
rect 24553 731 24583 783
rect 24447 729 24503 731
rect 24527 729 24583 731
rect 25271 783 25327 785
rect 25351 783 25407 785
rect 25271 731 25301 783
rect 25301 731 25313 783
rect 25313 731 25327 783
rect 25351 731 25365 783
rect 25365 731 25377 783
rect 25377 731 25407 783
rect 25271 729 25327 731
rect 25351 729 25407 731
rect 26051 783 26107 785
rect 26131 783 26187 785
rect 26051 731 26081 783
rect 26081 731 26093 783
rect 26093 731 26107 783
rect 26131 731 26145 783
rect 26145 731 26157 783
rect 26157 731 26187 783
rect 26051 729 26107 731
rect 26131 729 26187 731
rect 26831 783 26887 785
rect 26911 783 26967 785
rect 26831 731 26861 783
rect 26861 731 26873 783
rect 26873 731 26887 783
rect 26911 731 26925 783
rect 26925 731 26937 783
rect 26937 731 26967 783
rect 26831 729 26887 731
rect 26911 729 26967 731
<< metal3 >>
rect 200 7442 27389 7450
rect 200 7058 208 7442
rect 592 7058 12851 7442
rect 12995 7058 13675 7442
rect 13819 7058 14455 7442
rect 14599 7058 15235 7442
rect 15379 7058 24443 7442
rect 24587 7058 25267 7442
rect 25411 7058 26047 7442
rect 26191 7058 26827 7442
rect 26971 7058 27389 7442
rect 200 7052 27389 7058
rect 200 7050 600 7052
rect 12823 7050 13023 7052
rect 13647 7050 13847 7052
rect 14427 7050 14627 7052
rect 15207 7050 15407 7052
rect 24415 7050 24615 7052
rect 25239 7050 25439 7052
rect 26019 7050 26219 7052
rect 26799 7050 26999 7052
rect 200 6511 27389 6519
rect 200 6127 808 6511
rect 1192 6127 12458 6511
rect 12602 6127 13285 6511
rect 13429 6127 14065 6511
rect 14209 6127 14845 6511
rect 14989 6127 15625 6511
rect 15769 6127 24050 6511
rect 24194 6127 24877 6511
rect 25021 6127 25657 6511
rect 25801 6127 26437 6511
rect 26581 6127 27217 6511
rect 27361 6127 27389 6511
rect 200 6119 27389 6127
rect 12823 5501 13023 5509
rect 12823 5437 12851 5501
rect 12915 5437 12931 5501
rect 12995 5437 13023 5501
rect 12823 5429 13023 5437
rect 13647 5501 13847 5509
rect 13647 5437 13675 5501
rect 13739 5437 13755 5501
rect 13819 5437 13847 5501
rect 13647 5429 13847 5437
rect 14427 5501 14627 5509
rect 14427 5437 14455 5501
rect 14519 5437 14535 5501
rect 14599 5437 14627 5501
rect 14427 5429 14627 5437
rect 15207 5501 15407 5509
rect 15207 5437 15235 5501
rect 15299 5437 15315 5501
rect 15379 5437 15407 5501
rect 15207 5429 15407 5437
rect 24415 5501 24615 5509
rect 24415 5437 24443 5501
rect 24507 5437 24523 5501
rect 24587 5437 24615 5501
rect 24415 5429 24615 5437
rect 25239 5501 25439 5509
rect 25239 5437 25267 5501
rect 25331 5437 25347 5501
rect 25411 5437 25439 5501
rect 25239 5429 25439 5437
rect 26019 5501 26219 5509
rect 26019 5437 26047 5501
rect 26111 5437 26127 5501
rect 26191 5437 26219 5501
rect 26019 5429 26219 5437
rect 26799 5501 26999 5509
rect 26799 5437 26827 5501
rect 26891 5437 26907 5501
rect 26971 5437 26999 5501
rect 26799 5429 26999 5437
rect 12493 5364 15593 5369
rect 12493 5308 12502 5364
rect 12558 5308 13039 5364
rect 13095 5308 13329 5364
rect 13385 5308 13719 5364
rect 13775 5308 14109 5364
rect 14165 5308 14499 5364
rect 14555 5308 14889 5364
rect 14945 5308 15593 5364
rect 12493 5303 15593 5308
rect 24085 5364 27185 5369
rect 24085 5308 24094 5364
rect 24150 5308 24631 5364
rect 24687 5308 24921 5364
rect 24977 5308 25311 5364
rect 25367 5308 25701 5364
rect 25757 5308 26091 5364
rect 26147 5308 26481 5364
rect 26537 5308 27185 5364
rect 24085 5303 27185 5308
rect 13000 5095 15593 5113
rect 13000 5091 13675 5095
rect 13000 5035 13134 5091
rect 13190 5035 13394 5091
rect 13450 5035 13524 5091
rect 13580 5035 13675 5091
rect 13000 5031 13675 5035
rect 13739 5031 13755 5095
rect 13819 5091 14455 5095
rect 13840 5035 13914 5091
rect 13970 5035 14174 5091
rect 14230 5035 14304 5091
rect 14360 5035 14455 5091
rect 13819 5031 14455 5035
rect 14519 5031 14535 5095
rect 14599 5091 15235 5095
rect 14620 5035 14694 5091
rect 14750 5035 14954 5091
rect 15010 5035 15084 5091
rect 15140 5035 15235 5091
rect 14599 5031 15235 5035
rect 15299 5031 15315 5095
rect 15379 5031 15593 5095
rect 13000 5013 15593 5031
rect 24592 5095 27185 5113
rect 24592 5091 25267 5095
rect 24592 5035 24726 5091
rect 24782 5035 24986 5091
rect 25042 5035 25116 5091
rect 25172 5035 25267 5091
rect 24592 5031 25267 5035
rect 25331 5031 25347 5095
rect 25411 5091 26047 5095
rect 25432 5035 25506 5091
rect 25562 5035 25766 5091
rect 25822 5035 25896 5091
rect 25952 5035 26047 5091
rect 25411 5031 26047 5035
rect 26111 5031 26127 5095
rect 26191 5091 26827 5095
rect 26212 5035 26286 5091
rect 26342 5035 26546 5091
rect 26602 5035 26676 5091
rect 26732 5035 26827 5091
rect 26191 5031 26827 5035
rect 26891 5031 26907 5095
rect 26971 5031 27185 5095
rect 24592 5013 27185 5031
rect 15207 4930 15407 4931
rect 15207 4866 15235 4930
rect 15299 4866 15315 4930
rect 15379 4866 15407 4930
rect 15207 4865 15407 4866
rect 26799 4930 26999 4931
rect 26799 4866 26827 4930
rect 26891 4866 26907 4930
rect 26971 4866 26999 4930
rect 26799 4865 26999 4866
rect 15797 4301 18950 4302
rect 15797 4297 18788 4301
rect 15797 4241 15809 4297
rect 15865 4241 15889 4297
rect 15945 4241 18788 4297
rect 15797 4237 18788 4241
rect 18852 4237 18868 4301
rect 18932 4237 18950 4301
rect 15797 4236 18950 4237
rect 27389 4301 30542 4302
rect 27389 4297 30380 4301
rect 27389 4241 27401 4297
rect 27457 4241 27481 4297
rect 27537 4241 30380 4297
rect 27389 4237 30380 4241
rect 30444 4237 30460 4301
rect 30524 4237 30542 4301
rect 27389 4236 30542 4237
rect 15467 3594 15637 3595
rect 15467 3530 15480 3594
rect 15544 3530 15560 3594
rect 15624 3530 15637 3594
rect 15467 3529 15637 3530
rect 27059 3594 27229 3595
rect 27059 3530 27072 3594
rect 27136 3530 27152 3594
rect 27216 3530 27229 3594
rect 27059 3529 27229 3530
rect 12823 3451 15729 3469
rect 12823 3447 13285 3451
rect 11042 3404 12659 3405
rect 11042 3340 11060 3404
rect 11124 3340 11140 3404
rect 11204 3400 12659 3404
rect 11204 3344 12594 3400
rect 12650 3344 12659 3400
rect 12823 3391 13134 3447
rect 13190 3391 13285 3447
rect 12823 3387 13285 3391
rect 13349 3387 13365 3451
rect 13429 3447 14065 3451
rect 13450 3391 13524 3447
rect 13580 3391 13784 3447
rect 13840 3391 13914 3447
rect 13970 3391 14065 3447
rect 13429 3387 14065 3391
rect 14129 3387 14145 3451
rect 14209 3447 14845 3451
rect 14230 3391 14304 3447
rect 14360 3391 14564 3447
rect 14620 3391 14694 3447
rect 14750 3391 14845 3447
rect 14209 3387 14845 3391
rect 14909 3387 14925 3451
rect 14989 3447 15729 3451
rect 15010 3391 15084 3447
rect 15140 3391 15729 3447
rect 24415 3451 27321 3469
rect 24415 3447 24877 3451
rect 14989 3387 15729 3391
rect 12823 3369 15729 3387
rect 22634 3404 24251 3405
rect 11204 3340 12659 3344
rect 11042 3339 12659 3340
rect 22634 3340 22652 3404
rect 22716 3340 22732 3404
rect 22796 3400 24251 3404
rect 22796 3344 24186 3400
rect 24242 3344 24251 3400
rect 24415 3391 24726 3447
rect 24782 3391 24877 3447
rect 24415 3387 24877 3391
rect 24941 3387 24957 3451
rect 25021 3447 25657 3451
rect 25042 3391 25116 3447
rect 25172 3391 25376 3447
rect 25432 3391 25506 3447
rect 25562 3391 25657 3447
rect 25021 3387 25657 3391
rect 25721 3387 25737 3451
rect 25801 3447 26437 3451
rect 25822 3391 25896 3447
rect 25952 3391 26156 3447
rect 26212 3391 26286 3447
rect 26342 3391 26437 3447
rect 25801 3387 26437 3391
rect 26501 3387 26517 3451
rect 26581 3447 27321 3451
rect 26602 3391 26676 3447
rect 26732 3391 27321 3447
rect 26581 3387 27321 3391
rect 24415 3369 27321 3387
rect 22796 3340 24251 3344
rect 22634 3339 24251 3340
rect 12503 3274 16358 3279
rect 12503 3218 12686 3274
rect 12742 3218 13001 3274
rect 13057 3218 13329 3274
rect 13385 3218 13719 3274
rect 13775 3218 14109 3274
rect 14165 3218 14499 3274
rect 14555 3218 14889 3274
rect 14945 3265 16358 3274
rect 14945 3218 16196 3265
rect 12503 3213 16196 3218
rect 13257 3145 13457 3153
rect 13257 3081 13285 3145
rect 13349 3081 13365 3145
rect 13429 3081 13457 3145
rect 13257 3073 13457 3081
rect 14037 3145 14237 3153
rect 14037 3081 14065 3145
rect 14129 3081 14145 3145
rect 14209 3081 14237 3145
rect 14037 3073 14237 3081
rect 14817 3145 15017 3153
rect 14817 3081 14845 3145
rect 14909 3081 14925 3145
rect 14989 3081 15017 3145
rect 14817 3073 15017 3081
rect 16178 3013 16196 3213
rect 12677 3008 16196 3013
rect 12677 2952 12686 3008
rect 12742 2952 13329 3008
rect 13385 2952 13719 3008
rect 13775 2952 14109 3008
rect 14165 2952 14499 3008
rect 14555 2952 14889 3008
rect 14945 2952 15279 3008
rect 15335 2961 16196 3008
rect 16340 2961 16358 3265
rect 24095 3274 27950 3279
rect 24095 3218 24278 3274
rect 24334 3218 24593 3274
rect 24649 3218 24921 3274
rect 24977 3218 25311 3274
rect 25367 3218 25701 3274
rect 25757 3218 26091 3274
rect 26147 3218 26481 3274
rect 26537 3265 27950 3274
rect 26537 3218 27788 3265
rect 24095 3213 27788 3218
rect 24849 3145 25049 3153
rect 24849 3081 24877 3145
rect 24941 3081 24957 3145
rect 25021 3081 25049 3145
rect 24849 3073 25049 3081
rect 25629 3145 25829 3153
rect 25629 3081 25657 3145
rect 25721 3081 25737 3145
rect 25801 3081 25829 3145
rect 25629 3073 25829 3081
rect 26409 3145 26609 3153
rect 26409 3081 26437 3145
rect 26501 3081 26517 3145
rect 26581 3081 26609 3145
rect 26409 3073 26609 3081
rect 27770 3013 27788 3213
rect 15335 2952 16358 2961
rect 12677 2947 16358 2952
rect 24269 3008 27788 3013
rect 24269 2952 24278 3008
rect 24334 2952 24921 3008
rect 24977 2952 25311 3008
rect 25367 2952 25701 3008
rect 25757 2952 26091 3008
rect 26147 2952 26481 3008
rect 26537 2952 26871 3008
rect 26927 2961 27788 3008
rect 27932 2961 27950 3265
rect 26927 2952 27950 2961
rect 24269 2947 27950 2952
rect 13125 2839 15539 2857
rect 13125 2835 13285 2839
rect 13125 2779 13134 2835
rect 13190 2779 13264 2835
rect 13125 2775 13285 2779
rect 13349 2775 13365 2839
rect 13429 2835 14065 2839
rect 13429 2779 13524 2835
rect 13580 2779 13654 2835
rect 13710 2779 13914 2835
rect 13970 2779 14044 2835
rect 13429 2775 14065 2779
rect 14129 2775 14145 2839
rect 14209 2835 14845 2839
rect 14209 2779 14304 2835
rect 14360 2779 14434 2835
rect 14490 2779 14694 2835
rect 14750 2779 14824 2835
rect 14209 2775 14845 2779
rect 14909 2775 14925 2839
rect 14989 2835 15539 2839
rect 14989 2779 15084 2835
rect 15140 2779 15214 2835
rect 15270 2779 15474 2835
rect 15530 2779 15539 2835
rect 14989 2775 15539 2779
rect 13125 2757 15539 2775
rect 24717 2839 27131 2857
rect 24717 2835 24877 2839
rect 24717 2779 24726 2835
rect 24782 2779 24856 2835
rect 24717 2775 24877 2779
rect 24941 2775 24957 2839
rect 25021 2835 25657 2839
rect 25021 2779 25116 2835
rect 25172 2779 25246 2835
rect 25302 2779 25506 2835
rect 25562 2779 25636 2835
rect 25021 2775 25657 2779
rect 25721 2775 25737 2839
rect 25801 2835 26437 2839
rect 25801 2779 25896 2835
rect 25952 2779 26026 2835
rect 26082 2779 26286 2835
rect 26342 2779 26416 2835
rect 25801 2775 26437 2779
rect 26501 2775 26517 2839
rect 26581 2835 27131 2839
rect 26581 2779 26676 2835
rect 26732 2779 26806 2835
rect 26862 2779 27066 2835
rect 27122 2779 27131 2835
rect 26581 2775 27131 2779
rect 24717 2757 27131 2775
rect 12823 1195 15697 1213
rect 12823 1131 12851 1195
rect 12915 1131 12931 1195
rect 12995 1191 13675 1195
rect 12995 1135 13134 1191
rect 13190 1135 13264 1191
rect 13320 1135 13524 1191
rect 13580 1135 13654 1191
rect 12995 1131 13675 1135
rect 13739 1131 13755 1195
rect 13819 1191 14455 1195
rect 13819 1135 13914 1191
rect 13970 1135 14044 1191
rect 14100 1135 14304 1191
rect 14360 1135 14434 1191
rect 13819 1131 14455 1135
rect 14519 1131 14535 1195
rect 14599 1191 15235 1195
rect 14599 1135 14694 1191
rect 14750 1135 14824 1191
rect 14880 1135 15084 1191
rect 15140 1135 15214 1191
rect 14599 1131 15235 1135
rect 15299 1131 15315 1195
rect 15379 1191 15697 1195
rect 15379 1135 15474 1191
rect 15530 1135 15697 1191
rect 15379 1131 15697 1135
rect 12823 1113 15697 1131
rect 24415 1195 27289 1213
rect 24415 1131 24443 1195
rect 24507 1131 24523 1195
rect 24587 1191 25267 1195
rect 24587 1135 24726 1191
rect 24782 1135 24856 1191
rect 24912 1135 25116 1191
rect 25172 1135 25246 1191
rect 24587 1131 25267 1135
rect 25331 1131 25347 1195
rect 25411 1191 26047 1195
rect 25411 1135 25506 1191
rect 25562 1135 25636 1191
rect 25692 1135 25896 1191
rect 25952 1135 26026 1191
rect 25411 1131 26047 1135
rect 26111 1131 26127 1195
rect 26191 1191 26827 1195
rect 26191 1135 26286 1191
rect 26342 1135 26416 1191
rect 26472 1135 26676 1191
rect 26732 1135 26806 1191
rect 26191 1131 26827 1135
rect 26891 1131 26907 1195
rect 26971 1191 27289 1195
rect 26971 1135 27066 1191
rect 27122 1135 27289 1191
rect 26971 1131 27289 1135
rect 24415 1113 27289 1131
rect 12493 918 15697 923
rect 12493 862 12502 918
rect 12558 862 13329 918
rect 13385 862 13719 918
rect 13775 862 14109 918
rect 14165 862 14499 918
rect 14555 862 14889 918
rect 14945 862 15279 918
rect 15335 862 15697 918
rect 12493 857 15697 862
rect 24085 918 27289 923
rect 24085 862 24094 918
rect 24150 862 24921 918
rect 24977 862 25311 918
rect 25367 862 25701 918
rect 25757 862 26091 918
rect 26147 862 26481 918
rect 26537 862 26871 918
rect 26927 862 27289 918
rect 24085 857 27289 862
rect 12823 789 13023 797
rect 12823 725 12851 789
rect 12915 725 12931 789
rect 12995 725 13023 789
rect 12823 717 13023 725
rect 13647 789 13847 797
rect 13647 725 13675 789
rect 13739 725 13755 789
rect 13819 725 13847 789
rect 13647 717 13847 725
rect 14427 789 14627 797
rect 14427 725 14455 789
rect 14519 725 14535 789
rect 14599 725 14627 789
rect 14427 717 14627 725
rect 15207 789 15407 797
rect 15207 725 15235 789
rect 15299 725 15315 789
rect 15379 725 15407 789
rect 15207 717 15407 725
rect 24415 789 24615 797
rect 24415 725 24443 789
rect 24507 725 24523 789
rect 24587 725 24615 789
rect 24415 717 24615 725
rect 25239 789 25439 797
rect 25239 725 25267 789
rect 25331 725 25347 789
rect 25411 725 25439 789
rect 25239 717 25439 725
rect 26019 789 26219 797
rect 26019 725 26047 789
rect 26111 725 26127 789
rect 26191 725 26219 789
rect 26019 717 26219 725
rect 26799 789 26999 797
rect 26799 725 26827 789
rect 26891 725 26907 789
rect 26971 725 26999 789
rect 26799 717 26999 725
<< via3 >>
rect 208 7058 592 7442
rect 12851 7058 12995 7442
rect 13675 7058 13819 7442
rect 14455 7058 14599 7442
rect 15235 7058 15379 7442
rect 24443 7058 24587 7442
rect 25267 7058 25411 7442
rect 26047 7058 26191 7442
rect 26827 7058 26971 7442
rect 808 6127 1192 6511
rect 12458 6127 12602 6511
rect 13285 6127 13429 6511
rect 14065 6127 14209 6511
rect 14845 6127 14989 6511
rect 15625 6127 15769 6511
rect 24050 6127 24194 6511
rect 24877 6127 25021 6511
rect 25657 6127 25801 6511
rect 26437 6127 26581 6511
rect 27217 6127 27361 6511
rect 12851 5497 12915 5501
rect 12851 5441 12855 5497
rect 12855 5441 12911 5497
rect 12911 5441 12915 5497
rect 12851 5437 12915 5441
rect 12931 5497 12995 5501
rect 12931 5441 12935 5497
rect 12935 5441 12991 5497
rect 12991 5441 12995 5497
rect 12931 5437 12995 5441
rect 13675 5497 13739 5501
rect 13675 5441 13679 5497
rect 13679 5441 13735 5497
rect 13735 5441 13739 5497
rect 13675 5437 13739 5441
rect 13755 5497 13819 5501
rect 13755 5441 13759 5497
rect 13759 5441 13815 5497
rect 13815 5441 13819 5497
rect 13755 5437 13819 5441
rect 14455 5497 14519 5501
rect 14455 5441 14459 5497
rect 14459 5441 14515 5497
rect 14515 5441 14519 5497
rect 14455 5437 14519 5441
rect 14535 5497 14599 5501
rect 14535 5441 14539 5497
rect 14539 5441 14595 5497
rect 14595 5441 14599 5497
rect 14535 5437 14599 5441
rect 15235 5497 15299 5501
rect 15235 5441 15239 5497
rect 15239 5441 15295 5497
rect 15295 5441 15299 5497
rect 15235 5437 15299 5441
rect 15315 5497 15379 5501
rect 15315 5441 15319 5497
rect 15319 5441 15375 5497
rect 15375 5441 15379 5497
rect 15315 5437 15379 5441
rect 24443 5497 24507 5501
rect 24443 5441 24447 5497
rect 24447 5441 24503 5497
rect 24503 5441 24507 5497
rect 24443 5437 24507 5441
rect 24523 5497 24587 5501
rect 24523 5441 24527 5497
rect 24527 5441 24583 5497
rect 24583 5441 24587 5497
rect 24523 5437 24587 5441
rect 25267 5497 25331 5501
rect 25267 5441 25271 5497
rect 25271 5441 25327 5497
rect 25327 5441 25331 5497
rect 25267 5437 25331 5441
rect 25347 5497 25411 5501
rect 25347 5441 25351 5497
rect 25351 5441 25407 5497
rect 25407 5441 25411 5497
rect 25347 5437 25411 5441
rect 26047 5497 26111 5501
rect 26047 5441 26051 5497
rect 26051 5441 26107 5497
rect 26107 5441 26111 5497
rect 26047 5437 26111 5441
rect 26127 5497 26191 5501
rect 26127 5441 26131 5497
rect 26131 5441 26187 5497
rect 26187 5441 26191 5497
rect 26127 5437 26191 5441
rect 26827 5497 26891 5501
rect 26827 5441 26831 5497
rect 26831 5441 26887 5497
rect 26887 5441 26891 5497
rect 26827 5437 26891 5441
rect 26907 5497 26971 5501
rect 26907 5441 26911 5497
rect 26911 5441 26967 5497
rect 26967 5441 26971 5497
rect 26907 5437 26971 5441
rect 13675 5031 13739 5095
rect 13755 5091 13819 5095
rect 13755 5035 13784 5091
rect 13784 5035 13819 5091
rect 13755 5031 13819 5035
rect 14455 5031 14519 5095
rect 14535 5091 14599 5095
rect 14535 5035 14564 5091
rect 14564 5035 14599 5091
rect 14535 5031 14599 5035
rect 15235 5031 15299 5095
rect 15315 5031 15379 5095
rect 25267 5031 25331 5095
rect 25347 5091 25411 5095
rect 25347 5035 25376 5091
rect 25376 5035 25411 5091
rect 25347 5031 25411 5035
rect 26047 5031 26111 5095
rect 26127 5091 26191 5095
rect 26127 5035 26156 5091
rect 26156 5035 26191 5091
rect 26127 5031 26191 5035
rect 26827 5031 26891 5095
rect 26907 5031 26971 5095
rect 15235 4926 15299 4930
rect 15235 4870 15239 4926
rect 15239 4870 15295 4926
rect 15295 4870 15299 4926
rect 15235 4866 15299 4870
rect 15315 4926 15379 4930
rect 15315 4870 15319 4926
rect 15319 4870 15375 4926
rect 15375 4870 15379 4926
rect 15315 4866 15379 4870
rect 26827 4926 26891 4930
rect 26827 4870 26831 4926
rect 26831 4870 26887 4926
rect 26887 4870 26891 4926
rect 26827 4866 26891 4870
rect 26907 4926 26971 4930
rect 26907 4870 26911 4926
rect 26911 4870 26967 4926
rect 26967 4870 26971 4926
rect 26907 4866 26971 4870
rect 18788 4237 18852 4301
rect 18868 4237 18932 4301
rect 30380 4237 30444 4301
rect 30460 4237 30524 4301
rect 15480 3590 15544 3594
rect 15480 3534 15484 3590
rect 15484 3534 15540 3590
rect 15540 3534 15544 3590
rect 15480 3530 15544 3534
rect 15560 3590 15624 3594
rect 15560 3534 15564 3590
rect 15564 3534 15620 3590
rect 15620 3534 15624 3590
rect 15560 3530 15624 3534
rect 27072 3590 27136 3594
rect 27072 3534 27076 3590
rect 27076 3534 27132 3590
rect 27132 3534 27136 3590
rect 27072 3530 27136 3534
rect 27152 3590 27216 3594
rect 27152 3534 27156 3590
rect 27156 3534 27212 3590
rect 27212 3534 27216 3590
rect 27152 3530 27216 3534
rect 11060 3340 11124 3404
rect 11140 3340 11204 3404
rect 13285 3387 13349 3451
rect 13365 3447 13429 3451
rect 13365 3391 13394 3447
rect 13394 3391 13429 3447
rect 13365 3387 13429 3391
rect 14065 3387 14129 3451
rect 14145 3447 14209 3451
rect 14145 3391 14174 3447
rect 14174 3391 14209 3447
rect 14145 3387 14209 3391
rect 14845 3387 14909 3451
rect 14925 3447 14989 3451
rect 14925 3391 14954 3447
rect 14954 3391 14989 3447
rect 14925 3387 14989 3391
rect 22652 3340 22716 3404
rect 22732 3340 22796 3404
rect 24877 3387 24941 3451
rect 24957 3447 25021 3451
rect 24957 3391 24986 3447
rect 24986 3391 25021 3447
rect 24957 3387 25021 3391
rect 25657 3387 25721 3451
rect 25737 3447 25801 3451
rect 25737 3391 25766 3447
rect 25766 3391 25801 3447
rect 25737 3387 25801 3391
rect 26437 3387 26501 3451
rect 26517 3447 26581 3451
rect 26517 3391 26546 3447
rect 26546 3391 26581 3447
rect 26517 3387 26581 3391
rect 13285 3141 13349 3145
rect 13285 3085 13289 3141
rect 13289 3085 13345 3141
rect 13345 3085 13349 3141
rect 13285 3081 13349 3085
rect 13365 3141 13429 3145
rect 13365 3085 13369 3141
rect 13369 3085 13425 3141
rect 13425 3085 13429 3141
rect 13365 3081 13429 3085
rect 14065 3141 14129 3145
rect 14065 3085 14069 3141
rect 14069 3085 14125 3141
rect 14125 3085 14129 3141
rect 14065 3081 14129 3085
rect 14145 3141 14209 3145
rect 14145 3085 14149 3141
rect 14149 3085 14205 3141
rect 14205 3085 14209 3141
rect 14145 3081 14209 3085
rect 14845 3141 14909 3145
rect 14845 3085 14849 3141
rect 14849 3085 14905 3141
rect 14905 3085 14909 3141
rect 14845 3081 14909 3085
rect 14925 3141 14989 3145
rect 14925 3085 14929 3141
rect 14929 3085 14985 3141
rect 14985 3085 14989 3141
rect 14925 3081 14989 3085
rect 16196 2961 16340 3265
rect 24877 3141 24941 3145
rect 24877 3085 24881 3141
rect 24881 3085 24937 3141
rect 24937 3085 24941 3141
rect 24877 3081 24941 3085
rect 24957 3141 25021 3145
rect 24957 3085 24961 3141
rect 24961 3085 25017 3141
rect 25017 3085 25021 3141
rect 24957 3081 25021 3085
rect 25657 3141 25721 3145
rect 25657 3085 25661 3141
rect 25661 3085 25717 3141
rect 25717 3085 25721 3141
rect 25657 3081 25721 3085
rect 25737 3141 25801 3145
rect 25737 3085 25741 3141
rect 25741 3085 25797 3141
rect 25797 3085 25801 3141
rect 25737 3081 25801 3085
rect 26437 3141 26501 3145
rect 26437 3085 26441 3141
rect 26441 3085 26497 3141
rect 26497 3085 26501 3141
rect 26437 3081 26501 3085
rect 26517 3141 26581 3145
rect 26517 3085 26521 3141
rect 26521 3085 26577 3141
rect 26577 3085 26581 3141
rect 26517 3081 26581 3085
rect 27788 2961 27932 3265
rect 13285 2835 13349 2839
rect 13285 2779 13320 2835
rect 13320 2779 13349 2835
rect 13285 2775 13349 2779
rect 13365 2775 13429 2839
rect 14065 2835 14129 2839
rect 14065 2779 14100 2835
rect 14100 2779 14129 2835
rect 14065 2775 14129 2779
rect 14145 2775 14209 2839
rect 14845 2835 14909 2839
rect 14845 2779 14880 2835
rect 14880 2779 14909 2835
rect 14845 2775 14909 2779
rect 14925 2775 14989 2839
rect 24877 2835 24941 2839
rect 24877 2779 24912 2835
rect 24912 2779 24941 2835
rect 24877 2775 24941 2779
rect 24957 2775 25021 2839
rect 25657 2835 25721 2839
rect 25657 2779 25692 2835
rect 25692 2779 25721 2835
rect 25657 2775 25721 2779
rect 25737 2775 25801 2839
rect 26437 2835 26501 2839
rect 26437 2779 26472 2835
rect 26472 2779 26501 2835
rect 26437 2775 26501 2779
rect 26517 2775 26581 2839
rect 12851 1131 12915 1195
rect 12931 1131 12995 1195
rect 13675 1191 13739 1195
rect 13675 1135 13710 1191
rect 13710 1135 13739 1191
rect 13675 1131 13739 1135
rect 13755 1131 13819 1195
rect 14455 1191 14519 1195
rect 14455 1135 14490 1191
rect 14490 1135 14519 1191
rect 14455 1131 14519 1135
rect 14535 1131 14599 1195
rect 15235 1191 15299 1195
rect 15235 1135 15270 1191
rect 15270 1135 15299 1191
rect 15235 1131 15299 1135
rect 15315 1131 15379 1195
rect 24443 1131 24507 1195
rect 24523 1131 24587 1195
rect 25267 1191 25331 1195
rect 25267 1135 25302 1191
rect 25302 1135 25331 1191
rect 25267 1131 25331 1135
rect 25347 1131 25411 1195
rect 26047 1191 26111 1195
rect 26047 1135 26082 1191
rect 26082 1135 26111 1191
rect 26047 1131 26111 1135
rect 26127 1131 26191 1195
rect 26827 1191 26891 1195
rect 26827 1135 26862 1191
rect 26862 1135 26891 1191
rect 26827 1131 26891 1135
rect 26907 1131 26971 1195
rect 12851 785 12915 789
rect 12851 729 12855 785
rect 12855 729 12911 785
rect 12911 729 12915 785
rect 12851 725 12915 729
rect 12931 785 12995 789
rect 12931 729 12935 785
rect 12935 729 12991 785
rect 12991 729 12995 785
rect 12931 725 12995 729
rect 13675 785 13739 789
rect 13675 729 13679 785
rect 13679 729 13735 785
rect 13735 729 13739 785
rect 13675 725 13739 729
rect 13755 785 13819 789
rect 13755 729 13759 785
rect 13759 729 13815 785
rect 13815 729 13819 785
rect 13755 725 13819 729
rect 14455 785 14519 789
rect 14455 729 14459 785
rect 14459 729 14515 785
rect 14515 729 14519 785
rect 14455 725 14519 729
rect 14535 785 14599 789
rect 14535 729 14539 785
rect 14539 729 14595 785
rect 14595 729 14599 785
rect 14535 725 14599 729
rect 15235 785 15299 789
rect 15235 729 15239 785
rect 15239 729 15295 785
rect 15295 729 15299 785
rect 15235 725 15299 729
rect 15315 785 15379 789
rect 15315 729 15319 785
rect 15319 729 15375 785
rect 15375 729 15379 785
rect 15315 725 15379 729
rect 24443 785 24507 789
rect 24443 729 24447 785
rect 24447 729 24503 785
rect 24503 729 24507 785
rect 24443 725 24507 729
rect 24523 785 24587 789
rect 24523 729 24527 785
rect 24527 729 24583 785
rect 24583 729 24587 785
rect 24523 725 24587 729
rect 25267 785 25331 789
rect 25267 729 25271 785
rect 25271 729 25327 785
rect 25327 729 25331 785
rect 25267 725 25331 729
rect 25347 785 25411 789
rect 25347 729 25351 785
rect 25351 729 25407 785
rect 25407 729 25411 785
rect 25347 725 25411 729
rect 26047 785 26111 789
rect 26047 729 26051 785
rect 26051 729 26107 785
rect 26107 729 26111 785
rect 26047 725 26111 729
rect 26127 785 26191 789
rect 26127 729 26131 785
rect 26131 729 26187 785
rect 26187 729 26191 785
rect 26127 725 26191 729
rect 26827 785 26891 789
rect 26827 729 26831 785
rect 26831 729 26887 785
rect 26887 729 26891 785
rect 26827 725 26891 729
rect 26907 785 26971 789
rect 26907 729 26911 785
rect 26911 729 26967 785
rect 26967 729 26971 785
rect 26907 725 26971 729
<< metal4 >>
rect 6134 44152 6194 45152
rect 6686 44152 6746 45152
rect 7238 44152 7298 45152
rect 7790 44152 7850 45152
rect 8342 44152 8402 45152
rect 8894 44152 8954 45152
rect 9446 44152 9506 45152
rect 9998 44152 10058 45152
rect 10550 44152 10610 45152
rect 11102 44152 11162 45152
rect 11654 44152 11714 45152
rect 12206 44152 12266 45152
rect 12758 44152 12818 45152
rect 13310 44152 13370 45152
rect 13862 44152 13922 45152
rect 14414 44152 14474 45152
rect 14966 44152 15026 45152
rect 15518 44152 15578 45152
rect 16070 44152 16130 45152
rect 16622 44152 16682 45152
rect 17174 44152 17234 45152
rect 17726 44152 17786 45152
rect 18278 44152 18338 45152
rect 18830 44152 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 7442 600 44152
rect 200 7058 208 7442
rect 592 7058 600 7442
rect 200 1000 600 7058
rect 800 43952 18890 44152
rect 800 6511 1200 43952
rect 800 6127 808 6511
rect 1192 6127 1200 6511
rect 800 1000 1200 6127
rect 12430 6511 12630 7450
rect 12430 6127 12458 6511
rect 12602 6127 12630 6511
rect 11042 3404 11222 3405
rect 11042 3340 11060 3404
rect 11124 3340 11140 3404
rect 11204 3340 11222 3404
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 3340
rect 12430 717 12630 6127
rect 12823 7442 13023 7450
rect 12823 7058 12851 7442
rect 12995 7058 13023 7442
rect 12823 5501 13023 7058
rect 12823 5437 12851 5501
rect 12915 5437 12931 5501
rect 12995 5437 13023 5501
rect 12823 1195 13023 5437
rect 12823 1131 12851 1195
rect 12915 1131 12931 1195
rect 12995 1131 13023 1195
rect 12823 789 13023 1131
rect 12823 725 12851 789
rect 12915 725 12931 789
rect 12995 725 13023 789
rect 12823 717 13023 725
rect 13257 6511 13457 7450
rect 13257 6127 13285 6511
rect 13429 6127 13457 6511
rect 13257 3451 13457 6127
rect 13257 3387 13285 3451
rect 13349 3387 13365 3451
rect 13429 3387 13457 3451
rect 13257 3145 13457 3387
rect 13257 3081 13285 3145
rect 13349 3081 13365 3145
rect 13429 3081 13457 3145
rect 13257 2839 13457 3081
rect 13257 2775 13285 2839
rect 13349 2775 13365 2839
rect 13429 2775 13457 2839
rect 13257 717 13457 2775
rect 13647 7442 13847 7450
rect 13647 7058 13675 7442
rect 13819 7058 13847 7442
rect 13647 5501 13847 7058
rect 13647 5437 13675 5501
rect 13739 5437 13755 5501
rect 13819 5437 13847 5501
rect 13647 5095 13847 5437
rect 13647 5031 13675 5095
rect 13739 5031 13755 5095
rect 13819 5031 13847 5095
rect 13647 1195 13847 5031
rect 13647 1131 13675 1195
rect 13739 1131 13755 1195
rect 13819 1131 13847 1195
rect 13647 789 13847 1131
rect 13647 725 13675 789
rect 13739 725 13755 789
rect 13819 725 13847 789
rect 13647 717 13847 725
rect 14037 6511 14237 7450
rect 14037 6127 14065 6511
rect 14209 6127 14237 6511
rect 14037 3451 14237 6127
rect 14037 3387 14065 3451
rect 14129 3387 14145 3451
rect 14209 3387 14237 3451
rect 14037 3145 14237 3387
rect 14037 3081 14065 3145
rect 14129 3081 14145 3145
rect 14209 3081 14237 3145
rect 14037 2839 14237 3081
rect 14037 2775 14065 2839
rect 14129 2775 14145 2839
rect 14209 2775 14237 2839
rect 14037 717 14237 2775
rect 14427 7442 14627 7450
rect 14427 7058 14455 7442
rect 14599 7058 14627 7442
rect 14427 5501 14627 7058
rect 14427 5437 14455 5501
rect 14519 5437 14535 5501
rect 14599 5437 14627 5501
rect 14427 5095 14627 5437
rect 14427 5031 14455 5095
rect 14519 5031 14535 5095
rect 14599 5031 14627 5095
rect 14427 1195 14627 5031
rect 14427 1131 14455 1195
rect 14519 1131 14535 1195
rect 14599 1131 14627 1195
rect 14427 789 14627 1131
rect 14427 725 14455 789
rect 14519 725 14535 789
rect 14599 725 14627 789
rect 14427 717 14627 725
rect 14817 6511 15017 7450
rect 14817 6127 14845 6511
rect 14989 6127 15017 6511
rect 14817 3451 15017 6127
rect 14817 3387 14845 3451
rect 14909 3387 14925 3451
rect 14989 3387 15017 3451
rect 14817 3145 15017 3387
rect 14817 3081 14845 3145
rect 14909 3081 14925 3145
rect 14989 3081 15017 3145
rect 14817 2839 15017 3081
rect 14817 2775 14845 2839
rect 14909 2775 14925 2839
rect 14989 2775 15017 2839
rect 14817 717 15017 2775
rect 15207 7442 15407 7450
rect 15207 7058 15235 7442
rect 15379 7058 15407 7442
rect 15207 5501 15407 7058
rect 15207 5437 15235 5501
rect 15299 5437 15315 5501
rect 15379 5437 15407 5501
rect 15207 5095 15407 5437
rect 15207 5031 15235 5095
rect 15299 5031 15315 5095
rect 15379 5031 15407 5095
rect 15207 4930 15407 5031
rect 15207 4866 15235 4930
rect 15299 4866 15315 4930
rect 15379 4866 15407 4930
rect 15207 1195 15407 4866
rect 15597 6511 15797 7450
rect 15597 6127 15625 6511
rect 15769 6127 15797 6511
rect 15597 3595 15797 6127
rect 24022 6511 24222 7450
rect 24022 6127 24050 6511
rect 24194 6127 24222 6511
rect 15467 3594 15797 3595
rect 15467 3530 15480 3594
rect 15544 3530 15560 3594
rect 15624 3530 15797 3594
rect 15467 3529 15797 3530
rect 15207 1131 15235 1195
rect 15299 1131 15315 1195
rect 15379 1131 15407 1195
rect 15207 789 15407 1131
rect 15207 725 15235 789
rect 15299 725 15315 789
rect 15379 725 15407 789
rect 15207 717 15407 725
rect 15597 717 15797 3529
rect 18770 4301 18950 4302
rect 18770 4237 18788 4301
rect 18852 4237 18868 4301
rect 18932 4237 18950 4301
rect 16178 3265 16358 3279
rect 16178 2961 16196 3265
rect 16340 2961 16358 3265
rect 16178 480 16358 2961
rect 14906 300 16358 480
rect 14906 0 15086 300
rect 18770 0 18950 4237
rect 22634 3404 22814 3405
rect 22634 3340 22652 3404
rect 22716 3340 22732 3404
rect 22796 3340 22814 3404
rect 22634 0 22814 3340
rect 24022 717 24222 6127
rect 24415 7442 24615 7450
rect 24415 7058 24443 7442
rect 24587 7058 24615 7442
rect 24415 5501 24615 7058
rect 24415 5437 24443 5501
rect 24507 5437 24523 5501
rect 24587 5437 24615 5501
rect 24415 1195 24615 5437
rect 24415 1131 24443 1195
rect 24507 1131 24523 1195
rect 24587 1131 24615 1195
rect 24415 789 24615 1131
rect 24415 725 24443 789
rect 24507 725 24523 789
rect 24587 725 24615 789
rect 24415 717 24615 725
rect 24849 6511 25049 7450
rect 24849 6127 24877 6511
rect 25021 6127 25049 6511
rect 24849 3451 25049 6127
rect 24849 3387 24877 3451
rect 24941 3387 24957 3451
rect 25021 3387 25049 3451
rect 24849 3145 25049 3387
rect 24849 3081 24877 3145
rect 24941 3081 24957 3145
rect 25021 3081 25049 3145
rect 24849 2839 25049 3081
rect 24849 2775 24877 2839
rect 24941 2775 24957 2839
rect 25021 2775 25049 2839
rect 24849 717 25049 2775
rect 25239 7442 25439 7450
rect 25239 7058 25267 7442
rect 25411 7058 25439 7442
rect 25239 5501 25439 7058
rect 25239 5437 25267 5501
rect 25331 5437 25347 5501
rect 25411 5437 25439 5501
rect 25239 5095 25439 5437
rect 25239 5031 25267 5095
rect 25331 5031 25347 5095
rect 25411 5031 25439 5095
rect 25239 1195 25439 5031
rect 25239 1131 25267 1195
rect 25331 1131 25347 1195
rect 25411 1131 25439 1195
rect 25239 789 25439 1131
rect 25239 725 25267 789
rect 25331 725 25347 789
rect 25411 725 25439 789
rect 25239 717 25439 725
rect 25629 6511 25829 7450
rect 25629 6127 25657 6511
rect 25801 6127 25829 6511
rect 25629 3451 25829 6127
rect 25629 3387 25657 3451
rect 25721 3387 25737 3451
rect 25801 3387 25829 3451
rect 25629 3145 25829 3387
rect 25629 3081 25657 3145
rect 25721 3081 25737 3145
rect 25801 3081 25829 3145
rect 25629 2839 25829 3081
rect 25629 2775 25657 2839
rect 25721 2775 25737 2839
rect 25801 2775 25829 2839
rect 25629 717 25829 2775
rect 26019 7442 26219 7450
rect 26019 7058 26047 7442
rect 26191 7058 26219 7442
rect 26019 5501 26219 7058
rect 26019 5437 26047 5501
rect 26111 5437 26127 5501
rect 26191 5437 26219 5501
rect 26019 5095 26219 5437
rect 26019 5031 26047 5095
rect 26111 5031 26127 5095
rect 26191 5031 26219 5095
rect 26019 1195 26219 5031
rect 26019 1131 26047 1195
rect 26111 1131 26127 1195
rect 26191 1131 26219 1195
rect 26019 789 26219 1131
rect 26019 725 26047 789
rect 26111 725 26127 789
rect 26191 725 26219 789
rect 26019 717 26219 725
rect 26409 6511 26609 7450
rect 26409 6127 26437 6511
rect 26581 6127 26609 6511
rect 26409 3451 26609 6127
rect 26409 3387 26437 3451
rect 26501 3387 26517 3451
rect 26581 3387 26609 3451
rect 26409 3145 26609 3387
rect 26409 3081 26437 3145
rect 26501 3081 26517 3145
rect 26581 3081 26609 3145
rect 26409 2839 26609 3081
rect 26409 2775 26437 2839
rect 26501 2775 26517 2839
rect 26581 2775 26609 2839
rect 26409 717 26609 2775
rect 26799 7442 26999 7450
rect 26799 7058 26827 7442
rect 26971 7058 26999 7442
rect 26799 5501 26999 7058
rect 26799 5437 26827 5501
rect 26891 5437 26907 5501
rect 26971 5437 26999 5501
rect 26799 5095 26999 5437
rect 26799 5031 26827 5095
rect 26891 5031 26907 5095
rect 26971 5031 26999 5095
rect 26799 4930 26999 5031
rect 26799 4866 26827 4930
rect 26891 4866 26907 4930
rect 26971 4866 26999 4930
rect 26799 1195 26999 4866
rect 27189 6511 27389 7450
rect 27189 6127 27217 6511
rect 27361 6127 27389 6511
rect 27189 3595 27389 6127
rect 27059 3594 27389 3595
rect 27059 3530 27072 3594
rect 27136 3530 27152 3594
rect 27216 3530 27389 3594
rect 27059 3529 27389 3530
rect 26799 1131 26827 1195
rect 26891 1131 26907 1195
rect 26971 1131 26999 1195
rect 26799 789 26999 1131
rect 26799 725 26827 789
rect 26891 725 26907 789
rect 26971 725 26999 789
rect 26799 717 26999 725
rect 27189 717 27389 3529
rect 30362 4301 30542 4302
rect 30362 4237 30380 4301
rect 30444 4237 30460 4301
rect 30524 4237 30542 4301
rect 27770 3265 27950 3279
rect 27770 2961 27788 3265
rect 27932 2961 27950 3265
rect 27770 480 27950 2961
rect 26498 300 27950 480
rect 26498 0 26678 300
rect 30362 0 30542 4237
<< labels >>
flabel metal3 25486 5063 25486 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 25876 5063 25876 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 26266 5063 26266 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 24802 1163 24802 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 25192 1163 25192 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 25582 1163 25582 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 25972 1163 25972 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 26362 1163 26362 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 26752 1163 26752 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 26656 5063 26656 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 25096 5063 25096 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 25135 5336 25135 5336 2 FreeSans 480 0 0 0 vctrp
flabel metal3 13894 5063 13894 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 14284 5063 14284 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 14674 5063 14674 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 13210 1163 13210 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 13600 1163 13600 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 13990 1163 13990 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 14380 1163 14380 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 14770 1163 14770 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 15160 1163 15160 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 15064 5063 15064 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 13504 5063 13504 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 13543 5336 13543 5336 2 FreeSans 480 0 0 0 vctrp
flabel metal4 s 24122 5429 24122 5429 2 FreeSans 480 0 0 0 vss
flabel metal4 s 27289 5423 27289 5423 2 FreeSans 480 0 0 0 vss
flabel metal4 s 12530 5429 12530 5429 2 FreeSans 480 0 0 0 vss
flabel metal4 s 15697 5423 15697 5423 2 FreeSans 480 0 0 0 vss
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 600 90 0 0 clk
port 1 nsew
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 600 90 0 0 ena
port 2 nsew
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 600 90 0 0 rst_n
port 3 nsew
flabel metal4 s 30362 0 30542 200 0 FreeSans 1200 0 0 0 ua[0]
port 4 nsew
flabel metal4 s 26498 0 26678 200 0 FreeSans 1200 0 0 0 ua[1]
port 53 nsew
flabel metal4 s 22634 0 22814 200 0 FreeSans 1200 0 0 0 ua[2]
port 5 nsew
flabel metal4 s 18770 0 18950 200 0 FreeSans 1200 0 0 0 ua[3]
port 6 nsew
flabel metal4 s 14906 0 15086 200 0 FreeSans 1200 0 0 0 ua[4]
port 7 nsew
flabel metal4 s 11042 0 11222 200 0 FreeSans 1200 0 0 0 ua[5]
port 8 nsew
flabel metal4 s 7178 0 7358 200 0 FreeSans 1200 0 0 0 ua[6]
port 9 nsew
flabel metal4 s 3314 0 3494 200 0 FreeSans 1200 0 0 0 ua[7]
port 10 nsew
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 600 90 0 0 ui_in[0]
port 11 nsew
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 600 90 0 0 ui_in[1]
port 12 nsew
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 600 90 0 0 ui_in[2]
port 13 nsew
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 600 90 0 0 ui_in[3]
port 14 nsew
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 600 90 0 0 ui_in[4]
port 15 nsew
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 600 90 0 0 ui_in[5]
port 16 nsew
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 600 90 0 0 ui_in[6]
port 17 nsew
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 600 90 0 0 ui_in[7]
port 18 nsew
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 600 90 0 0 uio_in[0]
port 19 nsew
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 600 90 0 0 uio_in[1]
port 20 nsew
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 600 90 0 0 uio_in[2]
port 21 nsew
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 600 90 0 0 uio_in[3]
port 22 nsew
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 600 90 0 0 uio_in[4]
port 23 nsew
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 600 90 0 0 uio_in[5]
port 24 nsew
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 600 90 0 0 uio_in[6]
port 25 nsew
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 600 90 0 0 uio_in[7]
port 26 nsew
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 600 90 0 0 uio_oe[0]
port 27 nsew
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 600 90 0 0 uio_oe[1]
port 28 nsew
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 600 90 0 0 uio_oe[2]
port 29 nsew
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 600 90 0 0 uio_oe[3]
port 30 nsew
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 600 90 0 0 uio_oe[4]
port 31 nsew
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 600 90 0 0 uio_oe[5]
port 32 nsew
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 600 90 0 0 uio_oe[6]
port 33 nsew
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 600 90 0 0 uio_oe[7]
port 34 nsew
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 600 90 0 0 uio_out[0]
port 35 nsew
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 600 90 0 0 uio_out[1]
port 36 nsew
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 600 90 0 0 uio_out[2]
port 37 nsew
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 600 90 0 0 uio_out[3]
port 38 nsew
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 600 90 0 0 uio_out[4]
port 39 nsew
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 600 90 0 0 uio_out[5]
port 40 nsew
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 600 90 0 0 uio_out[6]
port 41 nsew
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 600 90 0 0 uio_out[7]
port 42 nsew
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 600 90 0 0 uo_out[0]
port 43 nsew
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 600 90 0 0 uo_out[1]
port 44 nsew
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 600 90 0 0 uo_out[2]
port 45 nsew
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 600 90 0 0 uo_out[3]
port 46 nsew
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 600 90 0 0 uo_out[4]
port 47 nsew
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 600 90 0 0 uo_out[5]
port 48 nsew
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 600 90 0 0 uo_out[6]
port 49 nsew
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 600 90 0 0 uo_out[7]
port 50 nsew
flabel metal4 s 200 1000 600 44152 1 FreeSans 500 0 0 0 VDPWR
port 51 nsew
flabel metal4 s 800 1000 1200 44152 1 FreeSans 500 0 0 0 VGND
port 52 nsew
flabel metal3 s 25207 5063 25207 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 s 25277 5336 25277 5336 2 FreeSans 480 0 0 0 vctrp
flabel metal3 s 25233 3419 25233 3419 2 FreeSans 480 0 0 0 vss
flabel metal3 s 25274 3246 25274 3246 2 FreeSans 480 0 0 0 vctrn
flabel metal3 s 25597 5063 25597 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 s 25667 5336 25667 5336 2 FreeSans 480 0 0 0 vctrp
flabel metal3 s 25623 3419 25623 3419 2 FreeSans 480 0 0 0 vss
flabel metal3 s 25664 3246 25664 3246 2 FreeSans 480 0 0 0 vctrn
flabel metal3 s 25987 5063 25987 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 s 26057 5336 26057 5336 2 FreeSans 480 0 0 0 vctrp
flabel metal3 s 26013 3419 26013 3419 2 FreeSans 480 0 0 0 vss
flabel metal3 s 26054 3246 26054 3246 2 FreeSans 480 0 0 0 vctrn
flabel metal3 s 25081 1163 25081 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 s 25011 890 25011 890 2 FreeSans 480 180 0 0 vctrp
flabel metal3 s 25055 2807 25055 2807 2 FreeSans 480 180 0 0 vss
flabel metal3 s 25014 2980 25014 2980 2 FreeSans 480 180 0 0 vctrn
flabel metal3 s 25471 1163 25471 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 s 25401 890 25401 890 2 FreeSans 480 180 0 0 vctrp
flabel metal3 s 25445 2807 25445 2807 2 FreeSans 480 180 0 0 vss
flabel metal3 s 25404 2980 25404 2980 2 FreeSans 480 180 0 0 vctrn
flabel metal3 s 25861 1163 25861 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 s 25791 890 25791 890 2 FreeSans 480 180 0 0 vctrp
flabel metal3 s 25835 2807 25835 2807 2 FreeSans 480 180 0 0 vss
flabel metal3 s 25794 2980 25794 2980 2 FreeSans 480 180 0 0 vctrn
flabel metal3 s 26251 1163 26251 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 s 26181 890 26181 890 2 FreeSans 480 180 0 0 vctrp
flabel metal3 s 26225 2807 26225 2807 2 FreeSans 480 180 0 0 vss
flabel metal3 s 26184 2980 26184 2980 2 FreeSans 480 180 0 0 vctrn
flabel metal3 s 26641 1163 26641 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 s 26571 890 26571 890 2 FreeSans 480 180 0 0 vctrp
flabel metal3 s 26615 2807 26615 2807 2 FreeSans 480 180 0 0 vss
flabel metal3 s 26574 2980 26574 2980 2 FreeSans 480 180 0 0 vctrn
flabel metal3 s 27031 1163 27031 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 s 26961 890 26961 890 2 FreeSans 480 180 0 0 vctrp
flabel metal3 s 27005 2807 27005 2807 2 FreeSans 480 180 0 0 vss
flabel metal3 s 26964 2980 26964 2980 2 FreeSans 480 180 0 0 vctrn
flabel metal3 s 26377 5063 26377 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 s 26447 5336 26447 5336 2 FreeSans 480 0 0 0 vctrp
flabel metal3 s 26403 3419 26403 3419 2 FreeSans 480 0 0 0 vss
flabel metal3 s 26444 3246 26444 3246 2 FreeSans 480 0 0 0 vctrn
flabel metal3 s 24817 5063 24817 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 s 24887 5336 24887 5336 2 FreeSans 480 0 0 0 vctrp
flabel metal3 s 24843 3419 24843 3419 2 FreeSans 480 0 0 0 vss
flabel metal3 s 24884 3246 24884 3246 2 FreeSans 480 0 0 0 vctrn
flabel metal3 s 24621 4737 24621 4737 2 FreeSans 480 0 0 0 vctrp
flabel metal3 s 24514 2980 24514 2980 2 FreeSans 480 0 0 0 vctrn
flabel metal3 s 24673 3419 24673 3419 2 FreeSans 480 0 0 0 vss
flabel metal3 s 24514 3246 24514 3246 2 FreeSans 480 0 0 0 vctrn
flabel metal3 s 24677 5063 24677 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 s 13615 5063 13615 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 s 13685 5336 13685 5336 2 FreeSans 480 0 0 0 vctrp
flabel metal3 s 13641 3419 13641 3419 2 FreeSans 480 0 0 0 vss
flabel metal3 s 13682 3246 13682 3246 2 FreeSans 480 0 0 0 vctrn
flabel metal3 s 14005 5063 14005 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 s 14075 5336 14075 5336 2 FreeSans 480 0 0 0 vctrp
flabel metal3 s 14031 3419 14031 3419 2 FreeSans 480 0 0 0 vss
flabel metal3 s 14072 3246 14072 3246 2 FreeSans 480 0 0 0 vctrn
flabel metal3 s 14395 5063 14395 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 s 14465 5336 14465 5336 2 FreeSans 480 0 0 0 vctrp
flabel metal3 s 14421 3419 14421 3419 2 FreeSans 480 0 0 0 vss
flabel metal3 s 14462 3246 14462 3246 2 FreeSans 480 0 0 0 vctrn
flabel metal3 s 13489 1163 13489 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 s 13419 890 13419 890 2 FreeSans 480 180 0 0 vctrp
flabel metal3 s 13463 2807 13463 2807 2 FreeSans 480 180 0 0 vss
flabel metal3 s 13422 2980 13422 2980 2 FreeSans 480 180 0 0 vctrn
flabel metal3 s 13879 1163 13879 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 s 13809 890 13809 890 2 FreeSans 480 180 0 0 vctrp
flabel metal3 s 13853 2807 13853 2807 2 FreeSans 480 180 0 0 vss
flabel metal3 s 13812 2980 13812 2980 2 FreeSans 480 180 0 0 vctrn
flabel metal3 s 14269 1163 14269 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 s 14199 890 14199 890 2 FreeSans 480 180 0 0 vctrp
flabel metal3 s 14243 2807 14243 2807 2 FreeSans 480 180 0 0 vss
flabel metal3 s 14202 2980 14202 2980 2 FreeSans 480 180 0 0 vctrn
flabel metal3 s 14659 1163 14659 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 s 14589 890 14589 890 2 FreeSans 480 180 0 0 vctrp
flabel metal3 s 14633 2807 14633 2807 2 FreeSans 480 180 0 0 vss
flabel metal3 s 14592 2980 14592 2980 2 FreeSans 480 180 0 0 vctrn
flabel metal3 s 15049 1163 15049 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 s 14979 890 14979 890 2 FreeSans 480 180 0 0 vctrp
flabel metal3 s 15023 2807 15023 2807 2 FreeSans 480 180 0 0 vss
flabel metal3 s 14982 2980 14982 2980 2 FreeSans 480 180 0 0 vctrn
flabel metal3 s 15439 1163 15439 1163 2 FreeSans 480 180 0 0 vdd
flabel metal3 s 15369 890 15369 890 2 FreeSans 480 180 0 0 vctrp
flabel metal3 s 15413 2807 15413 2807 2 FreeSans 480 180 0 0 vss
flabel metal3 s 15372 2980 15372 2980 2 FreeSans 480 180 0 0 vctrn
flabel metal3 s 14785 5063 14785 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 s 14855 5336 14855 5336 2 FreeSans 480 0 0 0 vctrp
flabel metal3 s 14811 3419 14811 3419 2 FreeSans 480 0 0 0 vss
flabel metal3 s 14852 3246 14852 3246 2 FreeSans 480 0 0 0 vctrn
flabel metal3 s 13225 5063 13225 5063 2 FreeSans 480 0 0 0 vdd
flabel metal3 s 13295 5336 13295 5336 2 FreeSans 480 0 0 0 vctrp
flabel metal3 s 13251 3419 13251 3419 2 FreeSans 480 0 0 0 vss
flabel metal3 s 13292 3246 13292 3246 2 FreeSans 480 0 0 0 vctrn
flabel metal3 s 13029 4737 13029 4737 2 FreeSans 480 0 0 0 vctrp
flabel metal3 s 12922 2980 12922 2980 2 FreeSans 480 0 0 0 vctrn
flabel metal3 s 13081 3419 13081 3419 2 FreeSans 480 0 0 0 vss
flabel metal3 s 12922 3246 12922 3246 2 FreeSans 480 0 0 0 vctrn
flabel metal3 s 13085 5063 13085 5063 2 FreeSans 480 0 0 0 vdd
flabel metal1 s 25154 4084 25154 4084 2 FreeSans 224 0 0 0 in
flabel metal1 s 25503 4086 25503 4086 2 FreeSans 224 0 0 0 out
flabel metal1 s 25302 5469 25302 5469 2 FreeSans 224 0 0 0 vdd
flabel metal1 s 25322 3112 25322 3112 2 FreeSans 224 0 0 0 vss
flabel metal1 s 25544 4084 25544 4084 2 FreeSans 224 0 0 0 in
flabel metal1 s 25893 4086 25893 4086 2 FreeSans 224 0 0 0 out
flabel metal1 s 25692 5469 25692 5469 2 FreeSans 224 0 0 0 vdd
flabel metal1 s 25712 3112 25712 3112 2 FreeSans 224 0 0 0 vss
flabel metal1 s 25934 4084 25934 4084 2 FreeSans 224 0 0 0 in
flabel metal1 s 26283 4086 26283 4086 2 FreeSans 224 0 0 0 out
flabel metal1 s 26082 5469 26082 5469 2 FreeSans 224 0 0 0 vdd
flabel metal1 s 26102 3112 26102 3112 2 FreeSans 224 0 0 0 vss
flabel metal1 s 25134 2142 25134 2142 2 FreeSans 224 180 0 0 in
flabel metal1 s 24785 2140 24785 2140 2 FreeSans 224 180 0 0 out
flabel metal1 s 24986 757 24986 757 2 FreeSans 224 180 0 0 vdd
flabel metal1 s 24966 3114 24966 3114 2 FreeSans 224 180 0 0 vss
flabel metal1 s 25524 2142 25524 2142 2 FreeSans 224 180 0 0 in
flabel metal1 s 25175 2140 25175 2140 2 FreeSans 224 180 0 0 out
flabel metal1 s 25376 757 25376 757 2 FreeSans 224 180 0 0 vdd
flabel metal1 s 25356 3114 25356 3114 2 FreeSans 224 180 0 0 vss
flabel metal1 s 25914 2142 25914 2142 2 FreeSans 224 180 0 0 in
flabel metal1 s 25565 2140 25565 2140 2 FreeSans 224 180 0 0 out
flabel metal1 s 25766 757 25766 757 2 FreeSans 224 180 0 0 vdd
flabel metal1 s 25746 3114 25746 3114 2 FreeSans 224 180 0 0 vss
flabel metal1 s 26304 2142 26304 2142 2 FreeSans 224 180 0 0 in
flabel metal1 s 25955 2140 25955 2140 2 FreeSans 224 180 0 0 out
flabel metal1 s 26156 757 26156 757 2 FreeSans 224 180 0 0 vdd
flabel metal1 s 26136 3114 26136 3114 2 FreeSans 224 180 0 0 vss
flabel metal1 s 26694 2142 26694 2142 2 FreeSans 224 180 0 0 in
flabel metal1 s 26345 2140 26345 2140 2 FreeSans 224 180 0 0 out
flabel metal1 s 26546 757 26546 757 2 FreeSans 224 180 0 0 vdd
flabel metal1 s 26526 3114 26526 3114 2 FreeSans 224 180 0 0 vss
flabel metal1 s 27084 2142 27084 2142 2 FreeSans 224 180 0 0 in
flabel metal1 s 26735 2140 26735 2140 2 FreeSans 224 180 0 0 out
flabel metal1 s 26936 757 26936 757 2 FreeSans 224 180 0 0 vdd
flabel metal1 s 26916 3114 26916 3114 2 FreeSans 224 180 0 0 vss
flabel metal1 s 26324 4084 26324 4084 2 FreeSans 224 0 0 0 in
flabel metal1 s 26673 4086 26673 4086 2 FreeSans 224 0 0 0 out
flabel metal1 s 26472 5469 26472 5469 2 FreeSans 224 0 0 0 vdd
flabel metal1 s 26492 3112 26492 3112 2 FreeSans 224 0 0 0 vss
flabel metal1 s 24764 4084 24764 4084 2 FreeSans 224 0 0 0 in
flabel metal1 s 25113 4086 25113 4086 2 FreeSans 224 0 0 0 out
flabel metal1 s 24912 5469 24912 5469 2 FreeSans 224 0 0 0 vdd
flabel metal1 s 24932 3112 24932 3112 2 FreeSans 224 0 0 0 vss
flabel metal1 s 27330 4279 27330 4279 2 FreeSans 224 0 0 0 out
flabel metal1 s 24528 3934 24528 3934 2 FreeSans 224 0 0 0 vrst
flabel metal1 s 24641 5469 24641 5469 2 FreeSans 224 0 0 0 vdd
flabel metal1 s 24597 3113 24597 3113 2 FreeSans 224 0 0 0 vss
flabel metal1 s 13562 4084 13562 4084 2 FreeSans 224 0 0 0 in
flabel metal1 s 13911 4086 13911 4086 2 FreeSans 224 0 0 0 out
flabel metal1 s 13710 5469 13710 5469 2 FreeSans 224 0 0 0 vdd
flabel metal1 s 13730 3112 13730 3112 2 FreeSans 224 0 0 0 vss
flabel metal1 s 13952 4084 13952 4084 2 FreeSans 224 0 0 0 in
flabel metal1 s 14301 4086 14301 4086 2 FreeSans 224 0 0 0 out
flabel metal1 s 14100 5469 14100 5469 2 FreeSans 224 0 0 0 vdd
flabel metal1 s 14120 3112 14120 3112 2 FreeSans 224 0 0 0 vss
flabel metal1 s 14342 4084 14342 4084 2 FreeSans 224 0 0 0 in
flabel metal1 s 14691 4086 14691 4086 2 FreeSans 224 0 0 0 out
flabel metal1 s 14490 5469 14490 5469 2 FreeSans 224 0 0 0 vdd
flabel metal1 s 14510 3112 14510 3112 2 FreeSans 224 0 0 0 vss
flabel metal1 s 13542 2142 13542 2142 2 FreeSans 224 180 0 0 in
flabel metal1 s 13193 2140 13193 2140 2 FreeSans 224 180 0 0 out
flabel metal1 s 13394 757 13394 757 2 FreeSans 224 180 0 0 vdd
flabel metal1 s 13374 3114 13374 3114 2 FreeSans 224 180 0 0 vss
flabel metal1 s 13932 2142 13932 2142 2 FreeSans 224 180 0 0 in
flabel metal1 s 13583 2140 13583 2140 2 FreeSans 224 180 0 0 out
flabel metal1 s 13784 757 13784 757 2 FreeSans 224 180 0 0 vdd
flabel metal1 s 13764 3114 13764 3114 2 FreeSans 224 180 0 0 vss
flabel metal1 s 14322 2142 14322 2142 2 FreeSans 224 180 0 0 in
flabel metal1 s 13973 2140 13973 2140 2 FreeSans 224 180 0 0 out
flabel metal1 s 14174 757 14174 757 2 FreeSans 224 180 0 0 vdd
flabel metal1 s 14154 3114 14154 3114 2 FreeSans 224 180 0 0 vss
flabel metal1 s 14712 2142 14712 2142 2 FreeSans 224 180 0 0 in
flabel metal1 s 14363 2140 14363 2140 2 FreeSans 224 180 0 0 out
flabel metal1 s 14564 757 14564 757 2 FreeSans 224 180 0 0 vdd
flabel metal1 s 14544 3114 14544 3114 2 FreeSans 224 180 0 0 vss
flabel metal1 s 15102 2142 15102 2142 2 FreeSans 224 180 0 0 in
flabel metal1 s 14753 2140 14753 2140 2 FreeSans 224 180 0 0 out
flabel metal1 s 14954 757 14954 757 2 FreeSans 224 180 0 0 vdd
flabel metal1 s 14934 3114 14934 3114 2 FreeSans 224 180 0 0 vss
flabel metal1 s 15492 2142 15492 2142 2 FreeSans 224 180 0 0 in
flabel metal1 s 15143 2140 15143 2140 2 FreeSans 224 180 0 0 out
flabel metal1 s 15344 757 15344 757 2 FreeSans 224 180 0 0 vdd
flabel metal1 s 15324 3114 15324 3114 2 FreeSans 224 180 0 0 vss
flabel metal1 s 14732 4084 14732 4084 2 FreeSans 224 0 0 0 in
flabel metal1 s 15081 4086 15081 4086 2 FreeSans 224 0 0 0 out
flabel metal1 s 14880 5469 14880 5469 2 FreeSans 224 0 0 0 vdd
flabel metal1 s 14900 3112 14900 3112 2 FreeSans 224 0 0 0 vss
flabel metal1 s 13172 4084 13172 4084 2 FreeSans 224 0 0 0 in
flabel metal1 s 13521 4086 13521 4086 2 FreeSans 224 0 0 0 out
flabel metal1 s 13320 5469 13320 5469 2 FreeSans 224 0 0 0 vdd
flabel metal1 s 13340 3112 13340 3112 2 FreeSans 224 0 0 0 vss
flabel metal1 s 15738 4279 15738 4279 2 FreeSans 224 0 0 0 out
flabel metal1 s 12936 3934 12936 3934 2 FreeSans 224 0 0 0 vrst
flabel metal1 s 13049 5469 13049 5469 2 FreeSans 224 0 0 0 vdd
flabel metal1 s 13005 3113 13005 3113 2 FreeSans 224 0 0 0 vss
<< properties >>
string FIXED_BBOX 0 0 32200 45152
string path 76.805 19.415 76.805 21.500 
<< end >>
